`timescale 1ns / 1ps

module streamGrp #(
    // hls4ml-streamGrp-gen-parameter
)(

    // hls4ml-streamGrp-gen-io

    input wire clk,
    input wire nreset

);

    // hls4ml-streamGrp-gen-create-module

endmodule