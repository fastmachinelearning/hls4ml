
//------> /opt/cad/catapult/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> /opt/cad/catapult/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  assign dat = idat;
  assign irdy = rdy;
  assign vld = ivld;

endmodule



//------> /opt/cad/catapult/pkgs/siflibs/ccs_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_vld_v1 (dat, vld, idat, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             vld;
  input  [width-1:0] idat;
  input              ivld;

  wire   [width-1:0] dat;
  wire               vld;

  assign dat = idat;
  assign vld = ivld;

endmodule


//------> /opt/cad/catapult/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/cad/catapult/pkgs/siflibs/mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ../td_ccore_solutions/nnet__sigmoid_layer4_t_result_t_sigmoid_config5__c9c110984abdfc2f0b91bec089345bc82281da_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4a/835166 Production Release
//  HLS Date:       Thu Sep  5 21:35:46 PDT 2019
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Mon Oct 21 13:59:08 2019
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    nnet_sigmoid_layer4_t_result_t_sigmoid_config5_core
// ------------------------------------------------------------------


module nnet_sigmoid_layer4_t_result_t_sigmoid_config5_core (
  data_rsc_dat, res_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_srst,
      ccs_ccore_en
);
  input [17:0] data_rsc_dat;
  output [17:0] res_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [17:0] data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg res_rsci_d_9;
  reg res_rsci_d_8;
  reg res_rsci_d_7;
  reg res_rsci_d_6;
  reg res_rsci_d_5;
  reg res_rsci_d_4;
  reg res_rsci_d_3;
  reg res_rsci_d_2;
  reg res_rsci_d_1;
  reg res_rsci_d_0;
  wire [5:0] index_14_9_lpi_1_dfm_1;
  wire sigmoid_table_and_cse;
  reg initialized_sva;
  reg sigmoid_table_511_2_sva;
  reg sigmoid_table_512_9_sva;
  reg sigmoid_table_510_3_sva;
  reg sigmoid_table_513_2_sva;
  reg sigmoid_table_513_9_sva;
  reg sigmoid_table_509_2_sva;
  reg sigmoid_table_509_4_sva;
  reg sigmoid_table_514_3_sva;
  reg sigmoid_table_514_9_sva;
  reg sigmoid_table_508_4_sva;
  reg sigmoid_table_515_2_sva;
  reg sigmoid_table_515_9_sva;
  reg sigmoid_table_507_2_sva;
  reg sigmoid_table_507_5_sva;
  reg sigmoid_table_516_0_sva;
  reg sigmoid_table_516_9_sva;
  reg sigmoid_table_506_3_sva;
  reg sigmoid_table_506_5_sva;
  reg sigmoid_table_517_4_sva;
  reg sigmoid_table_517_0_sva;
  reg sigmoid_table_517_9_sva;
  reg sigmoid_table_505_2_sva;
  reg sigmoid_table_505_5_sva;
  reg sigmoid_table_518_4_sva;
  reg sigmoid_table_518_0_sva;
  reg sigmoid_table_518_9_sva;
  reg sigmoid_table_504_5_sva;
  reg sigmoid_table_519_3_sva;
  reg sigmoid_table_519_0_sva;
  reg sigmoid_table_519_9_sva;
  reg sigmoid_table_503_2_sva;
  reg sigmoid_table_503_6_sva;
  reg sigmoid_table_520_0_sva;
  reg sigmoid_table_520_9_sva;
  reg sigmoid_table_502_3_sva;
  reg sigmoid_table_502_6_sva;
  reg sigmoid_table_521_5_sva;
  reg sigmoid_table_521_0_sva;
  reg sigmoid_table_521_9_sva;
  reg sigmoid_table_501_4_sva;
  reg sigmoid_table_501_2_sva;
  reg sigmoid_table_501_6_sva;
  reg sigmoid_table_522_5_sva;
  reg sigmoid_table_522_0_sva;
  reg sigmoid_table_522_9_sva;
  reg sigmoid_table_500_4_sva;
  reg sigmoid_table_500_6_sva;
  reg sigmoid_table_523_3_sva;
  reg sigmoid_table_523_5_sva;
  reg sigmoid_table_523_0_sva;
  reg sigmoid_table_523_9_sva;
  reg sigmoid_table_499_2_sva;
  reg sigmoid_table_499_6_sva;
  reg sigmoid_table_524_5_sva;
  reg sigmoid_table_524_0_sva;
  reg sigmoid_table_524_9_sva;
  reg sigmoid_table_498_3_sva;
  reg sigmoid_table_498_6_sva;
  reg sigmoid_table_525_4_sva;
  reg sigmoid_table_525_0_sva;
  reg sigmoid_table_525_9_sva;
  reg sigmoid_table_497_2_sva;
  reg sigmoid_table_497_6_sva;
  reg sigmoid_table_526_4_sva;
  reg sigmoid_table_526_0_sva;
  reg sigmoid_table_526_9_sva;
  reg sigmoid_table_496_6_sva;
  reg sigmoid_table_527_3_sva;
  reg sigmoid_table_527_0_sva;
  reg sigmoid_table_527_9_sva;
  reg sigmoid_table_495_2_sva;
  reg sigmoid_table_495_7_sva;
  reg sigmoid_table_528_0_sva;
  reg sigmoid_table_528_9_sva;
  reg sigmoid_table_494_3_sva;
  reg sigmoid_table_494_7_sva;
  reg sigmoid_table_529_6_sva;
  reg sigmoid_table_529_0_sva;
  reg sigmoid_table_529_9_sva;
  reg sigmoid_table_493_4_sva;
  reg sigmoid_table_493_2_sva;
  reg sigmoid_table_493_7_sva;
  reg sigmoid_table_530_6_sva;
  reg sigmoid_table_530_0_sva;
  reg sigmoid_table_530_9_sva;
  reg sigmoid_table_492_4_sva;
  reg sigmoid_table_492_7_sva;
  reg sigmoid_table_531_3_sva;
  reg sigmoid_table_531_6_sva;
  reg sigmoid_table_531_0_sva;
  reg sigmoid_table_531_9_sva;
  reg sigmoid_table_491_5_sva;
  reg sigmoid_table_491_2_sva;
  reg sigmoid_table_491_7_sva;
  reg sigmoid_table_532_6_sva;
  reg sigmoid_table_532_0_sva;
  reg sigmoid_table_532_9_sva;
  reg sigmoid_table_490_5_sva;
  reg sigmoid_table_490_3_sva;
  reg sigmoid_table_490_7_sva;
  reg sigmoid_table_533_4_sva;
  reg sigmoid_table_533_6_sva;
  reg sigmoid_table_533_0_sva;
  reg sigmoid_table_533_9_sva;
  reg sigmoid_table_489_5_sva;
  reg sigmoid_table_489_2_sva;
  reg sigmoid_table_489_7_sva;
  reg sigmoid_table_534_4_sva;
  reg sigmoid_table_534_6_sva;
  reg sigmoid_table_534_0_sva;
  reg sigmoid_table_534_9_sva;
  reg sigmoid_table_488_5_sva;
  reg sigmoid_table_488_0_sva;
  reg sigmoid_table_488_7_sva;
  reg sigmoid_table_535_3_sva;
  reg sigmoid_table_535_6_sva;
  reg sigmoid_table_535_0_sva;
  reg sigmoid_table_535_9_sva;
  reg sigmoid_table_487_2_sva;
  reg sigmoid_table_487_0_sva;
  reg sigmoid_table_487_7_sva;
  reg sigmoid_table_536_6_sva;
  reg sigmoid_table_536_1_sva;
  reg sigmoid_table_536_9_sva;
  reg sigmoid_table_486_3_sva;
  reg sigmoid_table_486_0_sva;
  reg sigmoid_table_486_7_sva;
  reg sigmoid_table_537_5_sva;
  reg sigmoid_table_537_1_sva;
  reg sigmoid_table_537_9_sva;
  reg sigmoid_table_485_2_sva;
  reg sigmoid_table_485_4_sva;
  reg sigmoid_table_485_0_sva;
  reg sigmoid_table_485_7_sva;
  reg sigmoid_table_538_5_sva;
  reg sigmoid_table_538_1_sva;
  reg sigmoid_table_538_9_sva;
  reg sigmoid_table_484_4_sva;
  reg sigmoid_table_484_0_sva;
  reg sigmoid_table_484_7_sva;
  reg sigmoid_table_539_3_sva;
  reg sigmoid_table_539_5_sva;
  reg sigmoid_table_539_1_sva;
  reg sigmoid_table_539_9_sva;
  reg sigmoid_table_483_2_sva;
  reg sigmoid_table_483_0_sva;
  reg sigmoid_table_483_7_sva;
  reg sigmoid_table_540_5_sva;
  reg sigmoid_table_540_1_sva;
  reg sigmoid_table_540_9_sva;
  reg sigmoid_table_482_3_sva;
  reg sigmoid_table_482_1_sva;
  reg sigmoid_table_482_7_sva;
  reg sigmoid_table_541_4_sva;
  reg sigmoid_table_541_1_sva;
  reg sigmoid_table_541_9_sva;
  reg sigmoid_table_481_1_sva;
  reg sigmoid_table_481_7_sva;
  reg sigmoid_table_542_2_sva;
  reg sigmoid_table_542_4_sva;
  reg sigmoid_table_542_0_sva;
  reg sigmoid_table_542_9_sva;
  reg sigmoid_table_480_1_sva;
  reg sigmoid_table_480_7_sva;
  reg sigmoid_table_543_3_sva;
  reg sigmoid_table_543_0_sva;
  reg sigmoid_table_543_9_sva;
  reg sigmoid_table_479_1_sva;
  reg sigmoid_table_479_8_sva;
  reg sigmoid_table_544_2_sva;
  reg sigmoid_table_544_0_sva;
  reg sigmoid_table_544_9_sva;
  reg sigmoid_table_478_3_sva;
  reg sigmoid_table_478_0_sva;
  reg sigmoid_table_478_8_sva;
  reg sigmoid_table_545_7_sva;
  reg sigmoid_table_545_0_sva;
  reg sigmoid_table_545_9_sva;
  reg sigmoid_table_477_4_sva;
  reg sigmoid_table_477_0_sva;
  reg sigmoid_table_477_8_sva;
  reg sigmoid_table_546_7_sva;
  reg sigmoid_table_546_2_sva;
  reg sigmoid_table_546_9_sva;
  reg sigmoid_table_476_4_sva;
  reg sigmoid_table_476_0_sva;
  reg sigmoid_table_476_8_sva;
  reg sigmoid_table_547_7_sva;
  reg sigmoid_table_547_3_sva;
  reg sigmoid_table_547_9_sva;
  reg sigmoid_table_475_5_sva;
  reg sigmoid_table_475_0_sva;
  reg sigmoid_table_475_8_sva;
  reg sigmoid_table_548_7_sva;
  reg sigmoid_table_548_2_sva;
  reg sigmoid_table_548_9_sva;
  reg sigmoid_table_474_5_sva;
  reg sigmoid_table_474_2_sva;
  reg sigmoid_table_474_8_sva;
  reg sigmoid_table_549_7_sva;
  reg sigmoid_table_549_4_sva;
  reg sigmoid_table_549_9_sva;
  reg sigmoid_table_473_5_sva;
  reg sigmoid_table_473_3_sva;
  reg sigmoid_table_473_8_sva;
  reg sigmoid_table_550_4_sva;
  reg sigmoid_table_550_7_sva;
  reg sigmoid_table_550_0_sva;
  reg sigmoid_table_550_9_sva;
  reg sigmoid_table_472_2_sva;
  reg sigmoid_table_472_5_sva;
  reg sigmoid_table_472_0_sva;
  reg sigmoid_table_472_8_sva;
  reg sigmoid_table_551_4_sva;
  reg sigmoid_table_551_7_sva;
  reg sigmoid_table_551_0_sva;
  reg sigmoid_table_551_9_sva;
  reg sigmoid_table_471_5_sva;
  reg sigmoid_table_471_0_sva;
  reg sigmoid_table_471_8_sva;
  reg sigmoid_table_552_3_sva;
  reg sigmoid_table_552_7_sva;
  reg sigmoid_table_552_1_sva;
  reg sigmoid_table_552_9_sva;
  reg sigmoid_table_470_2_sva;
  reg sigmoid_table_470_6_sva;
  reg sigmoid_table_470_0_sva;
  reg sigmoid_table_470_8_sva;
  reg sigmoid_table_553_7_sva;
  reg sigmoid_table_553_1_sva;
  reg sigmoid_table_553_9_sva;
  reg sigmoid_table_469_3_sva;
  reg sigmoid_table_469_6_sva;
  reg sigmoid_table_469_1_sva;
  reg sigmoid_table_469_8_sva;
  reg sigmoid_table_554_5_sva;
  reg sigmoid_table_554_7_sva;
  reg sigmoid_table_554_1_sva;
  reg sigmoid_table_554_9_sva;
  reg sigmoid_table_468_4_sva;
  reg sigmoid_table_468_6_sva;
  reg sigmoid_table_468_1_sva;
  reg sigmoid_table_468_8_sva;
  reg sigmoid_table_555_5_sva;
  reg sigmoid_table_555_2_sva;
  reg sigmoid_table_555_7_sva;
  reg sigmoid_table_555_0_sva;
  reg sigmoid_table_555_9_sva;
  reg sigmoid_table_467_4_sva;
  reg sigmoid_table_467_6_sva;
  reg sigmoid_table_467_0_sva;
  reg sigmoid_table_467_8_sva;
  reg sigmoid_table_556_5_sva;
  reg sigmoid_table_556_3_sva;
  reg sigmoid_table_556_7_sva;
  reg sigmoid_table_556_0_sva;
  reg sigmoid_table_556_9_sva;
  reg sigmoid_table_466_6_sva;
  reg sigmoid_table_466_0_sva;
  reg sigmoid_table_466_8_sva;
  reg sigmoid_table_557_5_sva;
  reg sigmoid_table_557_7_sva;
  reg sigmoid_table_557_2_sva;
  reg sigmoid_table_557_9_sva;
  reg sigmoid_table_465_6_sva;
  reg sigmoid_table_465_2_sva;
  reg sigmoid_table_465_8_sva;
  reg sigmoid_table_558_7_sva;
  reg sigmoid_table_558_4_sva;
  reg sigmoid_table_558_9_sva;
  reg sigmoid_table_464_6_sva;
  reg sigmoid_table_464_3_sva;
  reg sigmoid_table_464_8_sva;
  reg sigmoid_table_559_4_sva;
  reg sigmoid_table_559_7_sva;
  reg sigmoid_table_559_0_sva;
  reg sigmoid_table_559_9_sva;
  reg sigmoid_table_463_2_sva;
  reg sigmoid_table_463_6_sva;
  reg sigmoid_table_463_0_sva;
  reg sigmoid_table_463_8_sva;
  reg sigmoid_table_560_4_sva;
  reg sigmoid_table_560_7_sva;
  reg sigmoid_table_560_0_sva;
  reg sigmoid_table_560_9_sva;
  reg sigmoid_table_462_6_sva;
  reg sigmoid_table_462_0_sva;
  reg sigmoid_table_462_8_sva;
  reg sigmoid_table_561_3_sva;
  reg sigmoid_table_561_7_sva;
  reg sigmoid_table_561_1_sva;
  reg sigmoid_table_561_9_sva;
  reg sigmoid_table_461_1_sva;
  reg sigmoid_table_461_8_sva;
  reg sigmoid_table_562_7_sva;
  reg sigmoid_table_562_1_sva;
  reg sigmoid_table_562_9_sva;
  reg sigmoid_table_460_3_sva;
  reg sigmoid_table_460_1_sva;
  reg sigmoid_table_460_8_sva;
  reg sigmoid_table_563_6_sva;
  reg sigmoid_table_563_0_sva;
  reg sigmoid_table_563_9_sva;
  reg sigmoid_table_459_4_sva;
  reg sigmoid_table_459_0_sva;
  reg sigmoid_table_459_8_sva;
  reg sigmoid_table_564_2_sva;
  reg sigmoid_table_564_6_sva;
  reg sigmoid_table_564_0_sva;
  reg sigmoid_table_564_9_sva;
  reg sigmoid_table_458_4_sva;
  reg sigmoid_table_458_0_sva;
  reg sigmoid_table_458_8_sva;
  reg sigmoid_table_565_6_sva;
  reg sigmoid_table_565_3_sva;
  reg sigmoid_table_565_9_sva;
  reg sigmoid_table_457_4_sva;
  reg sigmoid_table_457_8_sva;
  reg sigmoid_table_566_6_sva;
  reg sigmoid_table_566_2_sva;
  reg sigmoid_table_566_9_sva;
  reg sigmoid_table_456_2_sva;
  reg sigmoid_table_456_5_sva;
  reg sigmoid_table_456_0_sva;
  reg sigmoid_table_456_8_sva;
  reg sigmoid_table_567_6_sva;
  reg sigmoid_table_567_0_sva;
  reg sigmoid_table_567_9_sva;
  reg sigmoid_table_455_3_sva;
  reg sigmoid_table_455_5_sva;
  reg sigmoid_table_455_0_sva;
  reg sigmoid_table_455_8_sva;
  reg sigmoid_table_568_4_sva;
  reg sigmoid_table_568_6_sva;
  reg sigmoid_table_568_1_sva;
  reg sigmoid_table_568_9_sva;
  reg sigmoid_table_454_5_sva;
  reg sigmoid_table_454_1_sva;
  reg sigmoid_table_454_8_sva;
  reg sigmoid_table_569_4_sva;
  reg sigmoid_table_569_6_sva;
  reg sigmoid_table_569_1_sva;
  reg sigmoid_table_569_9_sva;
  reg sigmoid_table_453_5_sva;
  reg sigmoid_table_453_0_sva;
  reg sigmoid_table_453_8_sva;
  reg sigmoid_table_570_3_sva;
  reg sigmoid_table_570_6_sva;
  reg sigmoid_table_570_0_sva;
  reg sigmoid_table_570_9_sva;
  reg sigmoid_table_452_5_sva;
  reg sigmoid_table_452_8_sva;
  reg sigmoid_table_571_6_sva;
  reg sigmoid_table_571_2_sva;
  reg sigmoid_table_571_9_sva;
  reg sigmoid_table_451_2_sva;
  reg sigmoid_table_451_8_sva;
  reg sigmoid_table_572_6_sva;
  reg sigmoid_table_572_0_sva;
  reg sigmoid_table_572_9_sva;
  reg sigmoid_table_450_3_sva;
  reg sigmoid_table_450_0_sva;
  reg sigmoid_table_450_8_sva;
  reg sigmoid_table_573_5_sva;
  reg sigmoid_table_573_0_sva;
  reg sigmoid_table_573_9_sva;
  reg sigmoid_table_449_4_sva;
  reg sigmoid_table_449_1_sva;
  reg sigmoid_table_449_8_sva;
  reg sigmoid_table_574_5_sva;
  reg sigmoid_table_574_1_sva;
  reg sigmoid_table_574_9_sva;
  reg sigmoid_table_448_4_sva;
  reg sigmoid_table_448_0_sva;
  reg sigmoid_table_448_8_sva;
  reg sigmoid_table_575_3_sva;
  reg sigmoid_table_575_5_sva;
  reg sigmoid_table_575_0_sva;
  reg sigmoid_table_575_9_sva;
  reg sigmoid_table_447_4_sva;
  reg sigmoid_table_447_8_sva;
  reg sigmoid_table_576_5_sva;
  reg sigmoid_table_576_2_sva;
  reg sigmoid_table_576_9_sva;
  reg sigmoid_table_446_2_sva;
  reg sigmoid_table_446_0_sva;
  reg sigmoid_table_446_8_sva;
  reg sigmoid_table_577_5_sva;
  reg sigmoid_table_577_0_sva;
  reg sigmoid_table_577_9_sva;
  reg sigmoid_table_445_3_sva;
  reg sigmoid_table_445_1_sva;
  reg sigmoid_table_445_8_sva;
  reg sigmoid_table_578_4_sva;
  reg sigmoid_table_578_1_sva;
  reg sigmoid_table_578_9_sva;
  reg sigmoid_table_444_1_sva;
  reg sigmoid_table_444_8_sva;
  reg sigmoid_table_579_2_sva;
  reg sigmoid_table_579_4_sva;
  reg sigmoid_table_579_0_sva;
  reg sigmoid_table_579_9_sva;
  reg sigmoid_table_443_0_sva;
  reg sigmoid_table_443_8_sva;
  reg sigmoid_table_580_3_sva;
  reg sigmoid_table_580_0_sva;
  reg sigmoid_table_580_9_sva;
  reg sigmoid_table_442_8_sva;
  reg sigmoid_table_581_2_sva;
  reg sigmoid_table_581_9_sva;
  reg sigmoid_table_441_0_sva;
  reg sigmoid_table_441_2_sva;
  reg sigmoid_table_582_0_sva;
  reg sigmoid_table_582_9_sva;
  reg sigmoid_table_440_1_sva;
  reg sigmoid_table_440_3_sva;
  reg sigmoid_table_583_1_sva;
  reg sigmoid_table_583_8_sva;
  reg sigmoid_table_439_3_sva;
  reg sigmoid_table_584_2_sva;
  reg sigmoid_table_584_0_sva;
  reg sigmoid_table_584_8_sva;
  reg sigmoid_table_438_2_sva;
  reg sigmoid_table_438_0_sva;
  reg sigmoid_table_438_4_sva;
  reg sigmoid_table_585_0_sva;
  reg sigmoid_table_585_8_sva;
  reg sigmoid_table_437_1_sva;
  reg sigmoid_table_437_4_sva;
  reg sigmoid_table_586_3_sva;
  reg sigmoid_table_586_1_sva;
  reg sigmoid_table_586_8_sva;
  reg sigmoid_table_436_0_sva;
  reg sigmoid_table_436_5_sva;
  reg sigmoid_table_587_2_sva;
  reg sigmoid_table_587_0_sva;
  reg sigmoid_table_587_8_sva;
  reg sigmoid_table_435_2_sva;
  reg sigmoid_table_435_5_sva;
  reg sigmoid_table_588_4_sva;
  reg sigmoid_table_588_8_sva;
  reg sigmoid_table_434_3_sva;
  reg sigmoid_table_434_0_sva;
  reg sigmoid_table_434_5_sva;
  reg sigmoid_table_589_4_sva;
  reg sigmoid_table_589_0_sva;
  reg sigmoid_table_589_8_sva;
  reg sigmoid_table_433_1_sva;
  reg sigmoid_table_433_5_sva;
  reg sigmoid_table_590_4_sva;
  reg sigmoid_table_590_1_sva;
  reg sigmoid_table_590_8_sva;
  reg sigmoid_table_432_2_sva;
  reg sigmoid_table_432_5_sva;
  reg sigmoid_table_591_3_sva;
  reg sigmoid_table_591_0_sva;
  reg sigmoid_table_591_8_sva;
  reg sigmoid_table_431_0_sva;
  reg sigmoid_table_431_5_sva;
  reg sigmoid_table_592_3_sva;
  reg sigmoid_table_592_0_sva;
  reg sigmoid_table_592_8_sva;
  reg sigmoid_table_430_1_sva;
  reg sigmoid_table_430_6_sva;
  reg sigmoid_table_593_1_sva;
  reg sigmoid_table_593_8_sva;
  reg sigmoid_table_429_3_sva;
  reg sigmoid_table_429_0_sva;
  reg sigmoid_table_429_6_sva;
  reg sigmoid_table_594_5_sva;
  reg sigmoid_table_594_0_sva;
  reg sigmoid_table_594_8_sva;
  reg sigmoid_table_428_3_sva;
  reg sigmoid_table_428_0_sva;
  reg sigmoid_table_428_6_sva;
  reg sigmoid_table_595_5_sva;
  reg sigmoid_table_595_2_sva;
  reg sigmoid_table_595_8_sva;
  reg sigmoid_table_427_4_sva;
  reg sigmoid_table_427_1_sva;
  reg sigmoid_table_427_6_sva;
  reg sigmoid_table_596_5_sva;
  reg sigmoid_table_596_1_sva;
  reg sigmoid_table_596_8_sva;
  reg sigmoid_table_426_4_sva;
  reg sigmoid_table_426_0_sva;
  reg sigmoid_table_426_6_sva;
  reg sigmoid_table_597_3_sva;
  reg sigmoid_table_597_5_sva;
  reg sigmoid_table_597_0_sva;
  reg sigmoid_table_597_8_sva;
  reg sigmoid_table_425_4_sva;
  reg sigmoid_table_425_0_sva;
  reg sigmoid_table_425_6_sva;
  reg sigmoid_table_598_5_sva;
  reg sigmoid_table_598_2_sva;
  reg sigmoid_table_598_8_sva;
  reg sigmoid_table_424_1_sva;
  reg sigmoid_table_424_6_sva;
  reg sigmoid_table_599_5_sva;
  reg sigmoid_table_599_1_sva;
  reg sigmoid_table_599_8_sva;
  reg sigmoid_table_423_2_sva;
  reg sigmoid_table_423_6_sva;
  reg sigmoid_table_600_4_sva;
  reg sigmoid_table_600_0_sva;
  reg sigmoid_table_600_8_sva;
  reg sigmoid_table_422_3_sva;
  reg sigmoid_table_422_0_sva;
  reg sigmoid_table_422_6_sva;
  reg sigmoid_table_601_4_sva;
  reg sigmoid_table_601_0_sva;
  reg sigmoid_table_601_8_sva;
  reg sigmoid_table_421_0_sva;
  reg sigmoid_table_421_6_sva;
  reg sigmoid_table_602_4_sva;
  reg sigmoid_table_602_1_sva;
  reg sigmoid_table_602_8_sva;
  reg sigmoid_table_420_2_sva;
  reg sigmoid_table_420_6_sva;
  reg sigmoid_table_603_3_sva;
  reg sigmoid_table_603_8_sva;
  reg sigmoid_table_419_1_sva;
  reg sigmoid_table_419_6_sva;
  reg sigmoid_table_604_3_sva;
  reg sigmoid_table_604_0_sva;
  reg sigmoid_table_604_8_sva;
  reg sigmoid_table_418_0_sva;
  reg sigmoid_table_418_7_sva;
  reg sigmoid_table_605_2_sva;
  reg sigmoid_table_605_0_sva;
  reg sigmoid_table_605_8_sva;
  reg sigmoid_table_417_2_sva;
  reg sigmoid_table_417_0_sva;
  reg sigmoid_table_417_7_sva;
  reg sigmoid_table_606_6_sva;
  reg sigmoid_table_606_8_sva;
  reg sigmoid_table_416_3_sva;
  reg sigmoid_table_416_1_sva;
  reg sigmoid_table_416_7_sva;
  reg sigmoid_table_607_6_sva;
  reg sigmoid_table_607_1_sva;
  reg sigmoid_table_607_8_sva;
  reg sigmoid_table_415_3_sva;
  reg sigmoid_table_415_7_sva;
  reg sigmoid_table_608_2_sva;
  reg sigmoid_table_608_6_sva;
  reg sigmoid_table_608_0_sva;
  reg sigmoid_table_608_8_sva;
  reg sigmoid_table_414_4_sva;
  reg sigmoid_table_414_1_sva;
  reg sigmoid_table_414_7_sva;
  reg sigmoid_table_609_6_sva;
  reg sigmoid_table_609_0_sva;
  reg sigmoid_table_609_8_sva;
  reg sigmoid_table_413_4_sva;
  reg sigmoid_table_413_0_sva;
  reg sigmoid_table_413_7_sva;
  reg sigmoid_table_610_3_sva;
  reg sigmoid_table_610_6_sva;
  reg sigmoid_table_610_0_sva;
  reg sigmoid_table_610_8_sva;
  reg sigmoid_table_412_4_sva;
  reg sigmoid_table_412_0_sva;
  reg sigmoid_table_412_7_sva;
  reg sigmoid_table_611_6_sva;
  reg sigmoid_table_611_2_sva;
  reg sigmoid_table_611_8_sva;
  reg sigmoid_table_411_5_sva;
  reg sigmoid_table_411_0_sva;
  reg sigmoid_table_411_7_sva;
  reg sigmoid_table_612_6_sva;
  reg sigmoid_table_612_1_sva;
  reg sigmoid_table_612_8_sva;
  reg sigmoid_table_410_5_sva;
  reg sigmoid_table_410_2_sva;
  reg sigmoid_table_410_7_sva;
  reg sigmoid_table_613_6_sva;
  reg sigmoid_table_613_4_sva;
  reg sigmoid_table_613_8_sva;
  reg sigmoid_table_409_3_sva;
  reg sigmoid_table_409_5_sva;
  reg sigmoid_table_409_1_sva;
  reg sigmoid_table_409_7_sva;
  reg sigmoid_table_614_4_sva;
  reg sigmoid_table_614_6_sva;
  reg sigmoid_table_614_0_sva;
  reg sigmoid_table_614_8_sva;
  reg sigmoid_table_408_5_sva;
  reg sigmoid_table_408_3_sva;
  reg sigmoid_table_408_7_sva;
  reg sigmoid_table_615_4_sva;
  reg sigmoid_table_615_2_sva;
  reg sigmoid_table_615_6_sva;
  reg sigmoid_table_615_0_sva;
  reg sigmoid_table_615_8_sva;
  reg sigmoid_table_407_5_sva;
  reg sigmoid_table_407_1_sva;
  reg sigmoid_table_407_7_sva;
  reg sigmoid_table_616_4_sva;
  reg sigmoid_table_616_6_sva;
  reg sigmoid_table_616_0_sva;
  reg sigmoid_table_616_8_sva;
  reg sigmoid_table_406_5_sva;
  reg sigmoid_table_406_2_sva;
  reg sigmoid_table_406_7_sva;
  reg sigmoid_table_617_3_sva;
  reg sigmoid_table_617_6_sva;
  reg sigmoid_table_617_0_sva;
  reg sigmoid_table_617_8_sva;
  reg sigmoid_table_405_5_sva;
  reg sigmoid_table_405_0_sva;
  reg sigmoid_table_405_7_sva;
  reg sigmoid_table_618_3_sva;
  reg sigmoid_table_618_6_sva;
  reg sigmoid_table_618_0_sva;
  reg sigmoid_table_618_8_sva;
  reg sigmoid_table_404_0_sva;
  reg sigmoid_table_404_7_sva;
  reg sigmoid_table_619_6_sva;
  reg sigmoid_table_619_1_sva;
  reg sigmoid_table_619_8_sva;
  reg sigmoid_table_403_2_sva;
  reg sigmoid_table_403_0_sva;
  reg sigmoid_table_403_7_sva;
  reg sigmoid_table_620_5_sva;
  reg sigmoid_table_620_8_sva;
  reg sigmoid_table_402_3_sva;
  reg sigmoid_table_402_0_sva;
  reg sigmoid_table_402_7_sva;
  reg sigmoid_table_621_5_sva;
  reg sigmoid_table_621_1_sva;
  reg sigmoid_table_621_8_sva;
  reg sigmoid_table_401_3_sva;
  reg sigmoid_table_401_0_sva;
  reg sigmoid_table_401_7_sva;
  reg sigmoid_table_622_5_sva;
  reg sigmoid_table_622_2_sva;
  reg sigmoid_table_622_8_sva;
  reg sigmoid_table_400_4_sva;
  reg sigmoid_table_400_0_sva;
  reg sigmoid_table_400_7_sva;
  reg sigmoid_table_623_5_sva;
  reg sigmoid_table_623_1_sva;
  reg sigmoid_table_623_8_sva;
  reg sigmoid_table_399_2_sva;
  reg sigmoid_table_399_4_sva;
  reg sigmoid_table_399_0_sva;
  reg sigmoid_table_399_7_sva;
  reg sigmoid_table_624_5_sva;
  reg sigmoid_table_624_3_sva;
  reg sigmoid_table_624_8_sva;
  reg sigmoid_table_398_4_sva;
  reg sigmoid_table_398_0_sva;
  reg sigmoid_table_398_7_sva;
  reg sigmoid_table_625_3_sva;
  reg sigmoid_table_625_5_sva;
  reg sigmoid_table_625_1_sva;
  reg sigmoid_table_625_8_sva;
  reg sigmoid_table_397_4_sva;
  reg sigmoid_table_397_0_sva;
  reg sigmoid_table_397_7_sva;
  reg sigmoid_table_626_5_sva;
  reg sigmoid_table_626_2_sva;
  reg sigmoid_table_626_8_sva;
  reg sigmoid_table_396_0_sva;
  reg sigmoid_table_396_7_sva;
  reg sigmoid_table_627_5_sva;
  reg sigmoid_table_627_1_sva;
  reg sigmoid_table_627_8_sva;
  reg sigmoid_table_395_2_sva;
  reg sigmoid_table_395_0_sva;
  reg sigmoid_table_395_7_sva;
  reg sigmoid_table_628_4_sva;
  reg sigmoid_table_628_8_sva;
  reg sigmoid_table_394_3_sva;
  reg sigmoid_table_394_0_sva;
  reg sigmoid_table_394_7_sva;
  reg sigmoid_table_629_4_sva;
  reg sigmoid_table_629_1_sva;
  reg sigmoid_table_629_8_sva;
  reg sigmoid_table_393_3_sva;
  reg sigmoid_table_393_1_sva;
  reg sigmoid_table_393_7_sva;
  reg sigmoid_table_630_4_sva;
  reg sigmoid_table_630_2_sva;
  reg sigmoid_table_630_8_sva;
  reg sigmoid_table_392_3_sva;
  reg sigmoid_table_392_7_sva;
  reg sigmoid_table_631_2_sva;
  reg sigmoid_table_631_4_sva;
  reg sigmoid_table_631_0_sva;
  reg sigmoid_table_631_8_sva;
  reg sigmoid_table_391_1_sva;
  reg sigmoid_table_391_7_sva;
  reg sigmoid_table_632_4_sva;
  reg sigmoid_table_632_0_sva;
  reg sigmoid_table_632_8_sva;
  reg sigmoid_table_390_2_sva;
  reg sigmoid_table_390_7_sva;
  reg sigmoid_table_633_3_sva;
  reg sigmoid_table_633_0_sva;
  reg sigmoid_table_633_8_sva;
  reg sigmoid_table_389_1_sva;
  reg sigmoid_table_389_7_sva;
  reg sigmoid_table_634_3_sva;
  reg sigmoid_table_634_0_sva;
  reg sigmoid_table_634_8_sva;
  reg sigmoid_table_388_7_sva;
  reg sigmoid_table_635_2_sva;
  reg sigmoid_table_635_0_sva;
  reg sigmoid_table_635_8_sva;
  reg sigmoid_table_387_0_sva;
  reg sigmoid_table_636_0_sva;
  reg sigmoid_table_636_8_sva;
  reg sigmoid_table_386_0_sva;
  reg sigmoid_table_386_2_sva;
  reg sigmoid_table_637_7_sva;
  reg sigmoid_table_385_0_sva;
  reg sigmoid_table_385_3_sva;
  reg sigmoid_table_638_1_sva;
  reg sigmoid_table_638_7_sva;
  reg sigmoid_table_384_1_sva;
  reg sigmoid_table_384_3_sva;
  reg sigmoid_table_639_2_sva;
  reg sigmoid_table_639_7_sva;
  reg sigmoid_table_383_3_sva;
  reg sigmoid_table_640_2_sva;
  reg sigmoid_table_640_0_sva;
  reg sigmoid_table_640_7_sva;
  reg sigmoid_table_382_1_sva;
  reg sigmoid_table_382_4_sva;
  reg sigmoid_table_641_0_sva;
  reg sigmoid_table_641_7_sva;
  reg sigmoid_table_381_2_sva;
  reg sigmoid_table_381_0_sva;
  reg sigmoid_table_381_4_sva;
  reg sigmoid_table_642_3_sva;
  reg sigmoid_table_642_0_sva;
  reg sigmoid_table_642_7_sva;
  reg sigmoid_table_380_0_sva;
  reg sigmoid_table_380_4_sva;
  reg sigmoid_table_643_3_sva;
  reg sigmoid_table_643_1_sva;
  reg sigmoid_table_643_7_sva;
  reg sigmoid_table_379_0_sva;
  reg sigmoid_table_379_4_sva;
  reg sigmoid_table_644_2_sva;
  reg sigmoid_table_644_7_sva;
  reg sigmoid_table_378_4_sva;
  reg sigmoid_table_645_1_sva;
  reg sigmoid_table_645_7_sva;
  reg sigmoid_table_377_1_sva;
  reg sigmoid_table_377_5_sva;
  reg sigmoid_table_646_0_sva;
  reg sigmoid_table_646_7_sva;
  reg sigmoid_table_376_2_sva;
  reg sigmoid_table_376_0_sva;
  reg sigmoid_table_376_5_sva;
  reg sigmoid_table_647_4_sva;
  reg sigmoid_table_647_0_sva;
  reg sigmoid_table_647_7_sva;
  reg sigmoid_table_375_3_sva;
  reg sigmoid_table_375_0_sva;
  reg sigmoid_table_375_5_sva;
  reg sigmoid_table_648_4_sva;
  reg sigmoid_table_648_1_sva;
  reg sigmoid_table_648_7_sva;
  reg sigmoid_table_374_3_sva;
  reg sigmoid_table_374_1_sva;
  reg sigmoid_table_374_5_sva;
  reg sigmoid_table_649_4_sva;
  reg sigmoid_table_649_2_sva;
  reg sigmoid_table_649_7_sva;
  reg sigmoid_table_373_3_sva;
  reg sigmoid_table_373_5_sva;
  reg sigmoid_table_650_2_sva;
  reg sigmoid_table_650_4_sva;
  reg sigmoid_table_650_0_sva;
  reg sigmoid_table_650_7_sva;
  reg sigmoid_table_372_0_sva;
  reg sigmoid_table_372_5_sva;
  reg sigmoid_table_651_4_sva;
  reg sigmoid_table_651_0_sva;
  reg sigmoid_table_651_7_sva;
  reg sigmoid_table_371_2_sva;
  reg sigmoid_table_371_0_sva;
  reg sigmoid_table_371_5_sva;
  reg sigmoid_table_652_3_sva;
  reg sigmoid_table_652_7_sva;
  reg sigmoid_table_370_2_sva;
  reg sigmoid_table_370_5_sva;
  reg sigmoid_table_653_3_sva;
  reg sigmoid_table_653_1_sva;
  reg sigmoid_table_653_7_sva;
  reg sigmoid_table_369_0_sva;
  reg sigmoid_table_369_5_sva;
  reg sigmoid_table_654_3_sva;
  reg sigmoid_table_654_0_sva;
  reg sigmoid_table_654_7_sva;
  reg sigmoid_table_368_0_sva;
  reg sigmoid_table_368_5_sva;
  reg sigmoid_table_655_2_sva;
  reg sigmoid_table_655_7_sva;
  reg sigmoid_table_367_5_sva;
  reg sigmoid_table_656_1_sva;
  reg sigmoid_table_656_7_sva;
  reg sigmoid_table_366_1_sva;
  reg sigmoid_table_366_6_sva;
  reg sigmoid_table_657_0_sva;
  reg sigmoid_table_657_7_sva;
  reg sigmoid_table_365_2_sva;
  reg sigmoid_table_365_0_sva;
  reg sigmoid_table_365_6_sva;
  reg sigmoid_table_658_5_sva;
  reg sigmoid_table_658_0_sva;
  reg sigmoid_table_658_7_sva;
  reg sigmoid_table_364_2_sva;
  reg sigmoid_table_364_6_sva;
  reg sigmoid_table_659_5_sva;
  reg sigmoid_table_659_1_sva;
  reg sigmoid_table_659_7_sva;
  reg sigmoid_table_363_3_sva;
  reg sigmoid_table_363_1_sva;
  reg sigmoid_table_363_6_sva;
  reg sigmoid_table_660_5_sva;
  reg sigmoid_table_660_0_sva;
  reg sigmoid_table_660_7_sva;
  reg sigmoid_table_362_3_sva;
  reg sigmoid_table_362_0_sva;
  reg sigmoid_table_362_6_sva;
  reg sigmoid_table_661_2_sva;
  reg sigmoid_table_661_5_sva;
  reg sigmoid_table_661_0_sva;
  reg sigmoid_table_661_7_sva;
  reg sigmoid_table_361_3_sva;
  reg sigmoid_table_361_6_sva;
  reg sigmoid_table_662_5_sva;
  reg sigmoid_table_662_1_sva;
  reg sigmoid_table_662_7_sva;
  reg sigmoid_table_360_4_sva;
  reg sigmoid_table_360_0_sva;
  reg sigmoid_table_360_6_sva;
  reg sigmoid_table_663_5_sva;
  reg sigmoid_table_663_0_sva;
  reg sigmoid_table_663_7_sva;
  reg sigmoid_table_359_2_sva;
  reg sigmoid_table_359_4_sva;
  reg sigmoid_table_359_0_sva;
  reg sigmoid_table_359_6_sva;
  reg sigmoid_table_664_5_sva;
  reg sigmoid_table_664_3_sva;
  reg sigmoid_table_664_7_sva;
  reg sigmoid_table_358_4_sva;
  reg sigmoid_table_358_2_sva;
  reg sigmoid_table_358_6_sva;
  reg sigmoid_table_665_3_sva;
  reg sigmoid_table_665_5_sva;
  reg sigmoid_table_665_1_sva;
  reg sigmoid_table_665_7_sva;
  reg sigmoid_table_357_4_sva;
  reg sigmoid_table_357_0_sva;
  reg sigmoid_table_357_6_sva;
  reg sigmoid_table_666_3_sva;
  reg sigmoid_table_666_5_sva;
  reg sigmoid_table_666_0_sva;
  reg sigmoid_table_666_7_sva;
  reg sigmoid_table_356_4_sva;
  reg sigmoid_table_356_1_sva;
  reg sigmoid_table_356_6_sva;
  reg sigmoid_table_667_5_sva;
  reg sigmoid_table_667_2_sva;
  reg sigmoid_table_667_7_sva;
  reg sigmoid_table_355_4_sva;
  reg sigmoid_table_355_0_sva;
  reg sigmoid_table_355_6_sva;
  reg sigmoid_table_668_2_sva;
  reg sigmoid_table_668_5_sva;
  reg sigmoid_table_668_0_sva;
  reg sigmoid_table_668_7_sva;
  reg sigmoid_table_354_0_sva;
  reg sigmoid_table_354_6_sva;
  reg sigmoid_table_669_5_sva;
  reg sigmoid_table_669_1_sva;
  reg sigmoid_table_669_7_sva;
  reg sigmoid_table_353_1_sva;
  reg sigmoid_table_353_6_sva;
  reg sigmoid_table_670_4_sva;
  reg sigmoid_table_670_7_sva;
  reg sigmoid_table_352_2_sva;
  reg sigmoid_table_352_0_sva;
  reg sigmoid_table_352_6_sva;
  reg sigmoid_table_671_4_sva;
  reg sigmoid_table_671_0_sva;
  reg sigmoid_table_671_7_sva;
  reg sigmoid_table_351_2_sva;
  reg sigmoid_table_351_6_sva;
  reg sigmoid_table_672_4_sva;
  reg sigmoid_table_672_1_sva;
  reg sigmoid_table_672_7_sva;
  reg sigmoid_table_350_3_sva;
  reg sigmoid_table_350_0_sva;
  reg sigmoid_table_350_6_sva;
  reg sigmoid_table_673_4_sva;
  reg sigmoid_table_673_0_sva;
  reg sigmoid_table_673_7_sva;
  reg sigmoid_table_349_3_sva;
  reg sigmoid_table_349_1_sva;
  reg sigmoid_table_349_6_sva;
  reg sigmoid_table_674_4_sva;
  reg sigmoid_table_674_2_sva;
  reg sigmoid_table_674_7_sva;
  reg sigmoid_table_348_3_sva;
  reg sigmoid_table_348_0_sva;
  reg sigmoid_table_348_6_sva;
  reg sigmoid_table_675_2_sva;
  reg sigmoid_table_675_4_sva;
  reg sigmoid_table_675_0_sva;
  reg sigmoid_table_675_7_sva;
  reg sigmoid_table_347_3_sva;
  reg sigmoid_table_347_6_sva;
  reg sigmoid_table_676_4_sva;
  reg sigmoid_table_676_1_sva;
  reg sigmoid_table_676_7_sva;
  reg sigmoid_table_346_0_sva;
  reg sigmoid_table_346_6_sva;
  reg sigmoid_table_677_4_sva;
  reg sigmoid_table_677_0_sva;
  reg sigmoid_table_677_7_sva;
  reg sigmoid_table_345_1_sva;
  reg sigmoid_table_345_6_sva;
  reg sigmoid_table_678_3_sva;
  reg sigmoid_table_678_7_sva;
  reg sigmoid_table_344_2_sva;
  reg sigmoid_table_344_0_sva;
  reg sigmoid_table_344_6_sva;
  reg sigmoid_table_679_3_sva;
  reg sigmoid_table_679_0_sva;
  reg sigmoid_table_679_7_sva;
  reg sigmoid_table_343_2_sva;
  reg sigmoid_table_343_6_sva;
  reg sigmoid_table_680_3_sva;
  reg sigmoid_table_680_1_sva;
  reg sigmoid_table_680_7_sva;
  reg sigmoid_table_342_0_sva;
  reg sigmoid_table_342_6_sva;
  reg sigmoid_table_681_3_sva;
  reg sigmoid_table_681_0_sva;
  reg sigmoid_table_681_7_sva;
  reg sigmoid_table_341_1_sva;
  reg sigmoid_table_341_6_sva;
  reg sigmoid_table_682_2_sva;
  reg sigmoid_table_682_7_sva;
  reg sigmoid_table_340_0_sva;
  reg sigmoid_table_340_6_sva;
  reg sigmoid_table_683_2_sva;
  reg sigmoid_table_683_0_sva;
  reg sigmoid_table_683_7_sva;
  reg sigmoid_table_339_6_sva;
  reg sigmoid_table_684_1_sva;
  reg sigmoid_table_684_7_sva;
  reg sigmoid_table_338_0_sva;
  reg sigmoid_table_685_0_sva;
  reg sigmoid_table_685_7_sva;
  reg sigmoid_table_337_1_sva;
  reg sigmoid_table_686_6_sva;
  reg sigmoid_table_336_0_sva;
  reg sigmoid_table_336_2_sva;
  reg sigmoid_table_687_0_sva;
  reg sigmoid_table_687_6_sva;
  reg sigmoid_table_335_2_sva;
  reg sigmoid_table_688_1_sva;
  reg sigmoid_table_688_6_sva;
  reg sigmoid_table_334_0_sva;
  reg sigmoid_table_334_3_sva;
  reg sigmoid_table_689_0_sva;
  reg sigmoid_table_689_6_sva;
  reg sigmoid_table_333_1_sva;
  reg sigmoid_table_333_3_sva;
  reg sigmoid_table_690_2_sva;
  reg sigmoid_table_690_6_sva;
  reg sigmoid_table_332_1_sva;
  reg sigmoid_table_332_3_sva;
  reg sigmoid_table_691_2_sva;
  reg sigmoid_table_691_0_sva;
  reg sigmoid_table_691_6_sva;
  reg sigmoid_table_331_0_sva;
  reg sigmoid_table_331_3_sva;
  reg sigmoid_table_692_2_sva;
  reg sigmoid_table_692_0_sva;
  reg sigmoid_table_692_6_sva;
  reg sigmoid_table_330_3_sva;
  reg sigmoid_table_693_1_sva;
  reg sigmoid_table_693_6_sva;
  reg sigmoid_table_329_0_sva;
  reg sigmoid_table_329_4_sva;
  reg sigmoid_table_694_0_sva;
  reg sigmoid_table_694_6_sva;
  reg sigmoid_table_328_1_sva;
  reg sigmoid_table_328_4_sva;
  reg sigmoid_table_695_3_sva;
  reg sigmoid_table_695_6_sva;
  reg sigmoid_table_327_2_sva;
  reg sigmoid_table_327_0_sva;
  reg sigmoid_table_327_4_sva;
  reg sigmoid_table_696_3_sva;
  reg sigmoid_table_696_0_sva;
  reg sigmoid_table_696_6_sva;
  reg sigmoid_table_326_2_sva;
  reg sigmoid_table_326_0_sva;
  reg sigmoid_table_326_4_sva;
  reg sigmoid_table_697_3_sva;
  reg sigmoid_table_697_1_sva;
  reg sigmoid_table_697_6_sva;
  reg sigmoid_table_325_2_sva;
  reg sigmoid_table_325_4_sva;
  reg sigmoid_table_698_3_sva;
  reg sigmoid_table_698_1_sva;
  reg sigmoid_table_698_6_sva;
  reg sigmoid_table_324_0_sva;
  reg sigmoid_table_324_4_sva;
  reg sigmoid_table_699_3_sva;
  reg sigmoid_table_699_0_sva;
  reg sigmoid_table_699_6_sva;
  reg sigmoid_table_323_1_sva;
  reg sigmoid_table_323_4_sva;
  reg sigmoid_table_700_2_sva;
  reg sigmoid_table_700_6_sva;
  reg sigmoid_table_322_1_sva;
  reg sigmoid_table_322_4_sva;
  reg sigmoid_table_701_2_sva;
  reg sigmoid_table_701_0_sva;
  reg sigmoid_table_701_6_sva;
  reg sigmoid_table_321_0_sva;
  reg sigmoid_table_321_4_sva;
  reg sigmoid_table_702_2_sva;
  reg sigmoid_table_702_0_sva;
  reg sigmoid_table_702_6_sva;
  reg sigmoid_table_320_4_sva;
  reg sigmoid_table_703_1_sva;
  reg sigmoid_table_703_6_sva;
  reg sigmoid_table_319_0_sva;
  reg sigmoid_table_319_5_sva;
  reg sigmoid_table_704_0_sva;
  reg sigmoid_table_704_6_sva;
  reg sigmoid_table_318_0_sva;
  reg sigmoid_table_318_5_sva;
  reg sigmoid_table_705_4_sva;
  reg sigmoid_table_705_6_sva;
  reg sigmoid_table_317_1_sva;
  reg sigmoid_table_317_5_sva;
  reg sigmoid_table_706_4_sva;
  reg sigmoid_table_706_6_sva;
  reg sigmoid_table_316_2_sva;
  reg sigmoid_table_316_0_sva;
  reg sigmoid_table_316_5_sva;
  reg sigmoid_table_707_4_sva;
  reg sigmoid_table_707_0_sva;
  reg sigmoid_table_707_6_sva;
  reg sigmoid_table_315_2_sva;
  reg sigmoid_table_315_0_sva;
  reg sigmoid_table_315_5_sva;
  reg sigmoid_table_708_4_sva;
  reg sigmoid_table_708_1_sva;
  reg sigmoid_table_708_6_sva;
  reg sigmoid_table_314_2_sva;
  reg sigmoid_table_314_5_sva;
  reg sigmoid_table_709_4_sva;
  reg sigmoid_table_709_1_sva;
  reg sigmoid_table_709_6_sva;
  reg sigmoid_table_313_3_sva;
  reg sigmoid_table_313_0_sva;
  reg sigmoid_table_313_5_sva;
  reg sigmoid_table_710_4_sva;
  reg sigmoid_table_710_0_sva;
  reg sigmoid_table_710_6_sva;
  reg sigmoid_table_312_3_sva;
  reg sigmoid_table_312_0_sva;
  reg sigmoid_table_312_5_sva;
  reg sigmoid_table_711_4_sva;
  reg sigmoid_table_711_2_sva;
  reg sigmoid_table_711_6_sva;
  reg sigmoid_table_311_3_sva;
  reg sigmoid_table_311_1_sva;
  reg sigmoid_table_311_5_sva;
  reg sigmoid_table_712_4_sva;
  reg sigmoid_table_712_2_sva;
  reg sigmoid_table_712_6_sva;
  reg sigmoid_table_310_3_sva;
  reg sigmoid_table_310_0_sva;
  reg sigmoid_table_310_5_sva;
  reg sigmoid_table_713_2_sva;
  reg sigmoid_table_713_4_sva;
  reg sigmoid_table_713_0_sva;
  reg sigmoid_table_713_6_sva;
  reg sigmoid_table_309_3_sva;
  reg sigmoid_table_309_0_sva;
  reg sigmoid_table_309_5_sva;
  reg sigmoid_table_714_4_sva;
  reg sigmoid_table_714_1_sva;
  reg sigmoid_table_714_6_sva;
  reg sigmoid_table_308_3_sva;
  reg sigmoid_table_308_5_sva;
  reg sigmoid_table_715_4_sva;
  reg sigmoid_table_715_1_sva;
  reg sigmoid_table_715_6_sva;
  reg sigmoid_table_307_0_sva;
  reg sigmoid_table_307_5_sva;
  reg sigmoid_table_716_4_sva;
  reg sigmoid_table_716_0_sva;
  reg sigmoid_table_716_6_sva;
  reg sigmoid_table_306_0_sva;
  reg sigmoid_table_306_5_sva;
  reg sigmoid_table_717_3_sva;
  reg sigmoid_table_717_6_sva;
  reg sigmoid_table_305_1_sva;
  reg sigmoid_table_305_5_sva;
  reg sigmoid_table_718_3_sva;
  reg sigmoid_table_718_6_sva;
  reg sigmoid_table_304_1_sva;
  reg sigmoid_table_304_5_sva;
  reg sigmoid_table_719_3_sva;
  reg sigmoid_table_719_0_sva;
  reg sigmoid_table_719_6_sva;
  reg sigmoid_table_303_2_sva;
  reg sigmoid_table_303_0_sva;
  reg sigmoid_table_303_5_sva;
  reg sigmoid_table_720_3_sva;
  reg sigmoid_table_720_0_sva;
  reg sigmoid_table_720_6_sva;
  reg sigmoid_table_302_2_sva;
  reg sigmoid_table_302_0_sva;
  reg sigmoid_table_302_5_sva;
  reg sigmoid_table_721_3_sva;
  reg sigmoid_table_721_1_sva;
  reg sigmoid_table_721_6_sva;
  reg sigmoid_table_301_2_sva;
  reg sigmoid_table_301_5_sva;
  reg sigmoid_table_722_3_sva;
  reg sigmoid_table_722_1_sva;
  reg sigmoid_table_722_6_sva;
  reg sigmoid_table_300_0_sva;
  reg sigmoid_table_300_5_sva;
  reg sigmoid_table_723_3_sva;
  reg sigmoid_table_723_0_sva;
  reg sigmoid_table_723_6_sva;
  reg sigmoid_table_299_0_sva;
  reg sigmoid_table_299_5_sva;
  reg sigmoid_table_724_2_sva;
  reg sigmoid_table_724_6_sva;
  reg sigmoid_table_298_1_sva;
  reg sigmoid_table_298_5_sva;
  reg sigmoid_table_725_2_sva;
  reg sigmoid_table_725_6_sva;
  reg sigmoid_table_297_1_sva;
  reg sigmoid_table_297_5_sva;
  reg sigmoid_table_726_2_sva;
  reg sigmoid_table_726_0_sva;
  reg sigmoid_table_726_6_sva;
  reg sigmoid_table_296_0_sva;
  reg sigmoid_table_296_5_sva;
  reg sigmoid_table_727_2_sva;
  reg sigmoid_table_727_0_sva;
  reg sigmoid_table_727_6_sva;
  reg sigmoid_table_295_0_sva;
  reg sigmoid_table_295_5_sva;
  reg sigmoid_table_728_1_sva;
  reg sigmoid_table_728_6_sva;
  reg sigmoid_table_294_5_sva;
  reg sigmoid_table_729_1_sva;
  reg sigmoid_table_729_6_sva;
  reg sigmoid_table_293_5_sva;
  reg sigmoid_table_730_0_sva;
  reg sigmoid_table_730_6_sva;
  reg sigmoid_table_292_0_sva;
  reg sigmoid_table_731_0_sva;
  reg sigmoid_table_731_6_sva;
  reg sigmoid_table_291_0_sva;
  reg sigmoid_table_732_5_sva;
  reg sigmoid_table_290_1_sva;
  reg sigmoid_table_733_5_sva;
  reg sigmoid_table_289_1_sva;
  reg sigmoid_table_734_0_sva;
  reg sigmoid_table_734_5_sva;
  reg sigmoid_table_288_1_sva;
  reg sigmoid_table_735_0_sva;
  reg sigmoid_table_735_5_sva;
  reg sigmoid_table_287_0_sva;
  reg sigmoid_table_287_2_sva;
  reg sigmoid_table_736_0_sva;
  reg sigmoid_table_736_5_sva;
  reg sigmoid_table_286_0_sva;
  reg sigmoid_table_286_2_sva;
  reg sigmoid_table_737_1_sva;
  reg sigmoid_table_737_5_sva;
  reg sigmoid_table_285_2_sva;
  reg sigmoid_table_738_1_sva;
  reg sigmoid_table_738_5_sva;
  reg sigmoid_table_284_2_sva;
  reg sigmoid_table_739_0_sva;
  reg sigmoid_table_739_5_sva;
  reg sigmoid_table_283_0_sva;
  reg sigmoid_table_283_3_sva;
  reg sigmoid_table_740_0_sva;
  reg sigmoid_table_740_5_sva;
  reg sigmoid_table_282_0_sva;
  reg sigmoid_table_282_3_sva;
  reg sigmoid_table_741_2_sva;
  reg sigmoid_table_741_5_sva;
  reg sigmoid_table_281_1_sva;
  reg sigmoid_table_281_3_sva;
  reg sigmoid_table_742_2_sva;
  reg sigmoid_table_742_5_sva;
  reg sigmoid_table_280_1_sva;
  reg sigmoid_table_280_3_sva;
  reg sigmoid_table_743_2_sva;
  reg sigmoid_table_743_0_sva;
  reg sigmoid_table_743_5_sva;
  reg sigmoid_table_279_1_sva;
  reg sigmoid_table_279_3_sva;
  reg sigmoid_table_744_2_sva;
  reg sigmoid_table_744_0_sva;
  reg sigmoid_table_744_5_sva;
  reg sigmoid_table_278_0_sva;
  reg sigmoid_table_278_3_sva;
  reg sigmoid_table_745_2_sva;
  reg sigmoid_table_745_0_sva;
  reg sigmoid_table_745_5_sva;
  reg sigmoid_table_277_0_sva;
  reg sigmoid_table_277_3_sva;
  reg sigmoid_table_746_1_sva;
  reg sigmoid_table_746_5_sva;
  reg sigmoid_table_276_0_sva;
  reg sigmoid_table_276_3_sva;
  reg sigmoid_table_747_1_sva;
  reg sigmoid_table_747_5_sva;
  reg sigmoid_table_275_3_sva;
  reg sigmoid_table_748_0_sva;
  reg sigmoid_table_748_5_sva;
  reg sigmoid_table_274_3_sva;
  reg sigmoid_table_749_0_sva;
  reg sigmoid_table_749_5_sva;
  reg sigmoid_table_273_0_sva;
  reg sigmoid_table_273_4_sva;
  reg sigmoid_table_750_0_sva;
  reg sigmoid_table_750_5_sva;
  reg sigmoid_table_272_0_sva;
  reg sigmoid_table_272_4_sva;
  reg sigmoid_table_751_3_sva;
  reg sigmoid_table_751_5_sva;
  reg sigmoid_table_271_0_sva;
  reg sigmoid_table_271_4_sva;
  reg sigmoid_table_752_3_sva;
  reg sigmoid_table_752_5_sva;
  reg sigmoid_table_270_1_sva;
  reg sigmoid_table_270_4_sva;
  reg sigmoid_table_753_3_sva;
  reg sigmoid_table_753_5_sva;
  reg sigmoid_table_269_1_sva;
  reg sigmoid_table_269_4_sva;
  reg sigmoid_table_754_3_sva;
  reg sigmoid_table_754_0_sva;
  reg sigmoid_table_754_5_sva;
  reg sigmoid_table_268_1_sva;
  reg sigmoid_table_268_4_sva;
  reg sigmoid_table_755_3_sva;
  reg sigmoid_table_755_0_sva;
  reg sigmoid_table_755_5_sva;
  reg sigmoid_table_267_2_sva;
  reg sigmoid_table_267_0_sva;
  reg sigmoid_table_267_4_sva;
  reg sigmoid_table_756_3_sva;
  reg sigmoid_table_756_0_sva;
  reg sigmoid_table_756_5_sva;
  reg sigmoid_table_266_2_sva;
  reg sigmoid_table_266_0_sva;
  reg sigmoid_table_266_4_sva;
  reg sigmoid_table_757_3_sva;
  reg sigmoid_table_757_1_sva;
  reg sigmoid_table_757_5_sva;
  reg sigmoid_table_265_2_sva;
  reg sigmoid_table_265_0_sva;
  reg sigmoid_table_265_4_sva;
  reg sigmoid_table_758_3_sva;
  reg sigmoid_table_758_1_sva;
  reg sigmoid_table_758_5_sva;
  reg sigmoid_table_264_2_sva;
  reg sigmoid_table_264_4_sva;
  reg sigmoid_table_759_3_sva;
  reg sigmoid_table_759_1_sva;
  reg sigmoid_table_759_5_sva;
  reg sigmoid_table_263_2_sva;
  reg sigmoid_table_263_4_sva;
  reg sigmoid_table_760_3_sva;
  reg sigmoid_table_760_0_sva;
  reg sigmoid_table_760_5_sva;
  reg sigmoid_table_262_2_sva;
  reg sigmoid_table_262_4_sva;
  reg sigmoid_table_761_3_sva;
  reg sigmoid_table_761_0_sva;
  reg sigmoid_table_761_5_sva;
  reg sigmoid_table_261_0_sva;
  reg sigmoid_table_261_4_sva;
  reg sigmoid_table_762_3_sva;
  reg sigmoid_table_762_0_sva;
  reg sigmoid_table_762_5_sva;
  reg sigmoid_table_260_0_sva;
  reg sigmoid_table_260_4_sva;
  reg sigmoid_table_763_2_sva;
  reg sigmoid_table_763_5_sva;
  reg sigmoid_table_259_0_sva;
  reg sigmoid_table_259_4_sva;
  reg sigmoid_table_764_2_sva;
  reg sigmoid_table_764_5_sva;
  reg sigmoid_table_258_1_sva;
  reg sigmoid_table_258_4_sva;
  reg sigmoid_table_765_2_sva;
  reg sigmoid_table_765_5_sva;
  reg sigmoid_table_257_1_sva;
  reg sigmoid_table_257_4_sva;
  reg sigmoid_table_766_2_sva;
  reg sigmoid_table_766_0_sva;
  reg sigmoid_table_766_5_sva;
  reg sigmoid_table_256_1_sva;
  reg sigmoid_table_256_4_sva;
  reg sigmoid_table_767_2_sva;
  reg sigmoid_table_767_0_sva;
  reg sigmoid_table_767_5_sva;
  reg sigmoid_table_255_1_sva;
  reg sigmoid_table_255_4_sva;
  reg sigmoid_table_768_2_sva;
  reg sigmoid_table_768_0_sva;
  reg sigmoid_table_768_5_sva;
  reg sigmoid_table_254_0_sva;
  reg sigmoid_table_254_4_sva;
  reg sigmoid_table_769_2_sva;
  reg sigmoid_table_769_0_sva;
  reg sigmoid_table_769_5_sva;
  reg sigmoid_table_253_0_sva;
  reg sigmoid_table_253_4_sva;
  reg sigmoid_table_770_1_sva;
  reg sigmoid_table_770_5_sva;
  reg sigmoid_table_252_0_sva;
  reg sigmoid_table_252_4_sva;
  reg sigmoid_table_771_1_sva;
  reg sigmoid_table_771_5_sva;
  reg sigmoid_table_251_0_sva;
  reg sigmoid_table_251_4_sva;
  reg sigmoid_table_772_1_sva;
  reg sigmoid_table_772_5_sva;
  reg sigmoid_table_250_4_sva;
  reg sigmoid_table_773_1_sva;
  reg sigmoid_table_773_5_sva;
  reg sigmoid_table_249_4_sva;
  reg sigmoid_table_774_0_sva;
  reg sigmoid_table_774_5_sva;
  reg sigmoid_table_248_4_sva;
  reg sigmoid_table_775_0_sva;
  reg sigmoid_table_775_5_sva;
  reg sigmoid_table_247_4_sva;
  reg sigmoid_table_776_0_sva;
  reg sigmoid_table_776_5_sva;
  reg sigmoid_table_246_0_sva;
  reg sigmoid_table_777_0_sva;
  reg sigmoid_table_777_5_sva;
  reg sigmoid_table_245_0_sva;
  reg sigmoid_table_778_4_sva;
  reg sigmoid_table_244_0_sva;
  reg sigmoid_table_779_4_sva;
  reg sigmoid_table_243_0_sva;
  reg sigmoid_table_780_4_sva;
  reg sigmoid_table_242_1_sva;
  reg sigmoid_table_781_4_sva;
  reg sigmoid_table_241_1_sva;
  reg sigmoid_table_782_0_sva;
  reg sigmoid_table_782_4_sva;
  reg sigmoid_table_240_1_sva;
  reg sigmoid_table_783_0_sva;
  reg sigmoid_table_783_4_sva;
  reg sigmoid_table_239_1_sva;
  reg sigmoid_table_784_0_sva;
  reg sigmoid_table_784_4_sva;
  reg sigmoid_table_238_0_sva;
  reg sigmoid_table_238_2_sva;
  reg sigmoid_table_785_0_sva;
  reg sigmoid_table_785_4_sva;
  reg sigmoid_table_237_0_sva;
  reg sigmoid_table_237_2_sva;
  reg sigmoid_table_786_1_sva;
  reg sigmoid_table_786_4_sva;
  reg sigmoid_table_236_0_sva;
  reg sigmoid_table_236_2_sva;
  reg sigmoid_table_787_1_sva;
  reg sigmoid_table_787_4_sva;
  reg sigmoid_table_235_0_sva;
  reg sigmoid_table_235_2_sva;
  reg sigmoid_table_788_1_sva;
  reg sigmoid_table_788_4_sva;
  reg sigmoid_table_234_0_sva;
  reg sigmoid_table_234_2_sva;
  reg sigmoid_table_789_1_sva;
  reg sigmoid_table_789_4_sva;
  reg sigmoid_table_233_2_sva;
  reg sigmoid_table_790_1_sva;
  reg sigmoid_table_790_4_sva;
  reg sigmoid_table_232_2_sva;
  reg sigmoid_table_791_0_sva;
  reg sigmoid_table_791_4_sva;
  reg sigmoid_table_231_2_sva;
  reg sigmoid_table_792_0_sva;
  reg sigmoid_table_792_4_sva;
  reg sigmoid_table_230_2_sva;
  reg sigmoid_table_793_0_sva;
  reg sigmoid_table_793_4_sva;
  reg sigmoid_table_229_2_sva;
  reg sigmoid_table_794_0_sva;
  reg sigmoid_table_794_4_sva;
  reg sigmoid_table_228_0_sva;
  reg sigmoid_table_228_3_sva;
  reg sigmoid_table_795_0_sva;
  reg sigmoid_table_795_4_sva;
  reg sigmoid_table_227_0_sva;
  reg sigmoid_table_227_3_sva;
  reg sigmoid_table_796_2_sva;
  reg sigmoid_table_796_4_sva;
  reg sigmoid_table_226_0_sva;
  reg sigmoid_table_226_3_sva;
  reg sigmoid_table_797_2_sva;
  reg sigmoid_table_797_4_sva;
  reg sigmoid_table_225_0_sva;
  reg sigmoid_table_225_3_sva;
  reg sigmoid_table_798_2_sva;
  reg sigmoid_table_798_4_sva;
  reg sigmoid_table_224_0_sva;
  reg sigmoid_table_224_3_sva;
  reg sigmoid_table_799_2_sva;
  reg sigmoid_table_799_4_sva;
  reg sigmoid_table_223_0_sva;
  reg sigmoid_table_223_3_sva;
  reg sigmoid_table_800_2_sva;
  reg sigmoid_table_800_4_sva;
  reg sigmoid_table_222_1_sva;
  reg sigmoid_table_222_3_sva;
  reg sigmoid_table_801_2_sva;
  reg sigmoid_table_801_4_sva;
  reg sigmoid_table_221_1_sva;
  reg sigmoid_table_221_3_sva;
  reg sigmoid_table_802_2_sva;
  reg sigmoid_table_802_0_sva;
  reg sigmoid_table_802_4_sva;
  reg sigmoid_table_220_1_sva;
  reg sigmoid_table_220_3_sva;
  reg sigmoid_table_803_2_sva;
  reg sigmoid_table_803_0_sva;
  reg sigmoid_table_803_4_sva;
  reg sigmoid_table_219_1_sva;
  reg sigmoid_table_219_3_sva;
  reg sigmoid_table_804_2_sva;
  reg sigmoid_table_804_0_sva;
  reg sigmoid_table_804_4_sva;
  reg sigmoid_table_218_1_sva;
  reg sigmoid_table_218_3_sva;
  reg sigmoid_table_805_2_sva;
  reg sigmoid_table_805_0_sva;
  reg sigmoid_table_805_4_sva;
  reg sigmoid_table_217_1_sva;
  reg sigmoid_table_217_3_sva;
  reg sigmoid_table_806_2_sva;
  reg sigmoid_table_806_0_sva;
  reg sigmoid_table_806_4_sva;
  reg sigmoid_table_216_0_sva;
  reg sigmoid_table_216_3_sva;
  reg sigmoid_table_807_2_sva;
  reg sigmoid_table_807_0_sva;
  reg sigmoid_table_807_4_sva;
  reg sigmoid_table_215_0_sva;
  reg sigmoid_table_215_3_sva;
  reg sigmoid_table_808_1_sva;
  reg sigmoid_table_808_4_sva;
  reg sigmoid_table_214_0_sva;
  reg sigmoid_table_214_3_sva;
  reg sigmoid_table_809_1_sva;
  reg sigmoid_table_809_4_sva;
  reg sigmoid_table_213_0_sva;
  reg sigmoid_table_213_3_sva;
  reg sigmoid_table_810_1_sva;
  reg sigmoid_table_810_4_sva;
  reg sigmoid_table_212_0_sva;
  reg sigmoid_table_212_3_sva;
  reg sigmoid_table_811_1_sva;
  reg sigmoid_table_811_4_sva;
  reg sigmoid_table_211_0_sva;
  reg sigmoid_table_211_3_sva;
  reg sigmoid_table_812_1_sva;
  reg sigmoid_table_812_4_sva;
  reg sigmoid_table_210_0_sva;
  reg sigmoid_table_210_3_sva;
  reg sigmoid_table_813_1_sva;
  reg sigmoid_table_813_4_sva;
  reg sigmoid_table_209_3_sva;
  reg sigmoid_table_814_1_sva;
  reg sigmoid_table_814_4_sva;
  reg sigmoid_table_208_3_sva;
  reg sigmoid_table_815_0_sva;
  reg sigmoid_table_815_4_sva;
  reg sigmoid_table_207_3_sva;
  reg sigmoid_table_816_0_sva;
  reg sigmoid_table_816_4_sva;
  reg sigmoid_table_206_3_sva;
  reg sigmoid_table_817_0_sva;
  reg sigmoid_table_817_4_sva;
  reg sigmoid_table_205_3_sva;
  reg sigmoid_table_818_0_sva;
  reg sigmoid_table_818_4_sva;
  reg sigmoid_table_204_3_sva;
  reg sigmoid_table_819_0_sva;
  reg sigmoid_table_819_4_sva;
  reg sigmoid_table_203_3_sva;
  reg sigmoid_table_820_0_sva;
  reg sigmoid_table_820_4_sva;
  reg sigmoid_table_202_3_sva;
  reg sigmoid_table_821_0_sva;
  reg sigmoid_table_821_4_sva;
  reg sigmoid_table_201_0_sva;
  reg sigmoid_table_822_3_sva;
  reg sigmoid_table_200_0_sva;
  reg sigmoid_table_823_3_sva;
  reg sigmoid_table_199_0_sva;
  reg sigmoid_table_824_3_sva;
  reg sigmoid_table_198_0_sva;
  reg sigmoid_table_825_3_sva;
  reg sigmoid_table_197_0_sva;
  reg sigmoid_table_826_3_sva;
  reg sigmoid_table_196_0_sva;
  reg sigmoid_table_827_3_sva;
  reg sigmoid_table_195_0_sva;
  reg sigmoid_table_828_3_sva;
  reg sigmoid_table_194_0_sva;
  reg sigmoid_table_829_3_sva;
  reg sigmoid_table_193_1_sva;
  reg sigmoid_table_830_3_sva;
  reg sigmoid_table_192_1_sva;
  reg sigmoid_table_831_0_sva;
  reg sigmoid_table_831_3_sva;
  reg sigmoid_table_191_1_sva;
  reg sigmoid_table_832_0_sva;
  reg sigmoid_table_832_3_sva;
  reg sigmoid_table_190_1_sva;
  reg sigmoid_table_833_0_sva;
  reg sigmoid_table_833_3_sva;
  reg sigmoid_table_189_1_sva;
  reg sigmoid_table_834_0_sva;
  reg sigmoid_table_834_3_sva;
  reg sigmoid_table_188_1_sva;
  reg sigmoid_table_835_0_sva;
  reg sigmoid_table_835_3_sva;
  reg sigmoid_table_187_1_sva;
  reg sigmoid_table_836_0_sva;
  reg sigmoid_table_836_3_sva;
  reg sigmoid_table_186_1_sva;
  reg sigmoid_table_837_0_sva;
  reg sigmoid_table_837_3_sva;
  reg sigmoid_table_185_1_sva;
  reg sigmoid_table_838_0_sva;
  reg sigmoid_table_838_3_sva;
  reg sigmoid_table_184_1_sva;
  reg sigmoid_table_839_0_sva;
  reg sigmoid_table_839_3_sva;
  reg sigmoid_table_183_0_sva;
  reg sigmoid_table_183_2_sva;
  reg sigmoid_table_840_0_sva;
  reg sigmoid_table_840_3_sva;
  reg sigmoid_table_182_0_sva;
  reg sigmoid_table_182_2_sva;
  reg sigmoid_table_841_1_sva;
  reg sigmoid_table_841_3_sva;
  reg sigmoid_table_181_0_sva;
  reg sigmoid_table_181_2_sva;
  reg sigmoid_table_842_1_sva;
  reg sigmoid_table_842_3_sva;
  reg sigmoid_table_180_0_sva;
  reg sigmoid_table_180_2_sva;
  reg sigmoid_table_843_1_sva;
  reg sigmoid_table_843_3_sva;
  reg sigmoid_table_179_0_sva;
  reg sigmoid_table_179_2_sva;
  reg sigmoid_table_844_1_sva;
  reg sigmoid_table_844_3_sva;
  reg sigmoid_table_178_0_sva;
  reg sigmoid_table_178_2_sva;
  reg sigmoid_table_845_1_sva;
  reg sigmoid_table_845_3_sva;
  reg sigmoid_table_177_0_sva;
  reg sigmoid_table_177_2_sva;
  reg sigmoid_table_846_1_sva;
  reg sigmoid_table_846_3_sva;
  reg sigmoid_table_176_0_sva;
  reg sigmoid_table_176_2_sva;
  reg sigmoid_table_847_1_sva;
  reg sigmoid_table_847_3_sva;
  reg sigmoid_table_175_0_sva;
  reg sigmoid_table_175_2_sva;
  reg sigmoid_table_848_1_sva;
  reg sigmoid_table_848_3_sva;
  reg sigmoid_table_174_0_sva;
  reg sigmoid_table_174_2_sva;
  reg sigmoid_table_849_1_sva;
  reg sigmoid_table_849_3_sva;
  reg sigmoid_table_173_0_sva;
  reg sigmoid_table_173_2_sva;
  reg sigmoid_table_850_1_sva;
  reg sigmoid_table_850_3_sva;
  reg sigmoid_table_172_0_sva;
  reg sigmoid_table_172_2_sva;
  reg sigmoid_table_851_1_sva;
  reg sigmoid_table_851_3_sva;
  reg sigmoid_table_171_2_sva;
  reg sigmoid_table_852_1_sva;
  reg sigmoid_table_852_3_sva;
  reg sigmoid_table_170_2_sva;
  reg sigmoid_table_853_0_sva;
  reg sigmoid_table_853_3_sva;
  reg sigmoid_table_169_2_sva;
  reg sigmoid_table_854_0_sva;
  reg sigmoid_table_854_3_sva;
  reg sigmoid_table_168_2_sva;
  reg sigmoid_table_855_0_sva;
  reg sigmoid_table_855_3_sva;
  reg sigmoid_table_167_2_sva;
  reg sigmoid_table_856_0_sva;
  reg sigmoid_table_856_3_sva;
  reg sigmoid_table_166_2_sva;
  reg sigmoid_table_857_0_sva;
  reg sigmoid_table_857_3_sva;
  reg sigmoid_table_165_2_sva;
  reg sigmoid_table_858_0_sva;
  reg sigmoid_table_858_3_sva;
  reg sigmoid_table_164_2_sva;
  reg sigmoid_table_859_0_sva;
  reg sigmoid_table_859_3_sva;
  reg sigmoid_table_163_2_sva;
  reg sigmoid_table_860_0_sva;
  reg sigmoid_table_860_3_sva;
  reg sigmoid_table_162_2_sva;
  reg sigmoid_table_861_0_sva;
  reg sigmoid_table_861_3_sva;
  reg sigmoid_table_161_2_sva;
  reg sigmoid_table_862_0_sva;
  reg sigmoid_table_862_3_sva;
  reg sigmoid_table_160_2_sva;
  reg sigmoid_table_863_0_sva;
  reg sigmoid_table_863_3_sva;
  reg sigmoid_table_159_2_sva;
  reg sigmoid_table_864_0_sva;
  reg sigmoid_table_864_3_sva;
  reg sigmoid_table_158_2_sva;
  reg sigmoid_table_865_0_sva;
  reg sigmoid_table_865_3_sva;
  reg sigmoid_table_157_0_sva;
  reg sigmoid_table_866_0_sva;
  reg sigmoid_table_866_3_sva;
  reg sigmoid_table_156_0_sva;
  reg sigmoid_table_867_2_sva;
  reg sigmoid_table_155_0_sva;
  reg sigmoid_table_868_2_sva;
  reg sigmoid_table_154_0_sva;
  reg sigmoid_table_869_2_sva;
  reg sigmoid_table_153_0_sva;
  reg sigmoid_table_870_2_sva;
  reg sigmoid_table_152_0_sva;
  reg sigmoid_table_871_2_sva;
  reg sigmoid_table_151_0_sva;
  reg sigmoid_table_872_2_sva;
  reg sigmoid_table_150_0_sva;
  reg sigmoid_table_873_2_sva;
  reg sigmoid_table_149_0_sva;
  reg sigmoid_table_874_2_sva;
  reg sigmoid_table_148_0_sva;
  reg sigmoid_table_875_2_sva;
  reg sigmoid_table_147_0_sva;
  reg sigmoid_table_876_2_sva;
  reg sigmoid_table_146_0_sva;
  reg sigmoid_table_877_2_sva;
  reg sigmoid_table_145_0_sva;
  reg sigmoid_table_878_2_sva;
  reg sigmoid_table_144_0_sva;
  reg sigmoid_table_879_2_sva;
  reg sigmoid_table_143_0_sva;
  reg sigmoid_table_880_2_sva;
  reg sigmoid_table_142_0_sva;
  reg sigmoid_table_881_2_sva;
  reg sigmoid_table_141_0_sva;
  reg sigmoid_table_882_2_sva;
  reg sigmoid_table_140_0_sva;
  reg sigmoid_table_883_2_sva;
  reg sigmoid_table_139_0_sva;
  reg sigmoid_table_884_2_sva;
  reg sigmoid_table_138_1_sva;
  reg sigmoid_table_885_0_sva;
  reg sigmoid_table_885_2_sva;
  reg sigmoid_table_137_1_sva;
  reg sigmoid_table_886_0_sva;
  reg sigmoid_table_886_2_sva;
  reg sigmoid_table_136_1_sva;
  reg sigmoid_table_887_0_sva;
  reg sigmoid_table_887_2_sva;
  reg sigmoid_table_135_1_sva;
  reg sigmoid_table_888_0_sva;
  reg sigmoid_table_888_2_sva;
  reg sigmoid_table_134_1_sva;
  reg sigmoid_table_889_0_sva;
  reg sigmoid_table_889_2_sva;
  reg sigmoid_table_133_1_sva;
  reg sigmoid_table_890_0_sva;
  reg sigmoid_table_890_2_sva;
  reg sigmoid_table_132_1_sva;
  reg sigmoid_table_891_0_sva;
  reg sigmoid_table_891_2_sva;
  reg sigmoid_table_131_1_sva;
  reg sigmoid_table_892_0_sva;
  reg sigmoid_table_892_2_sva;
  reg sigmoid_table_130_1_sva;
  reg sigmoid_table_893_0_sva;
  reg sigmoid_table_893_2_sva;
  reg sigmoid_table_129_1_sva;
  reg sigmoid_table_894_0_sva;
  reg sigmoid_table_894_2_sva;
  reg sigmoid_table_128_1_sva;
  reg sigmoid_table_895_0_sva;
  reg sigmoid_table_895_2_sva;
  reg sigmoid_table_127_1_sva;
  reg sigmoid_table_896_0_sva;
  reg sigmoid_table_896_2_sva;
  reg sigmoid_table_126_1_sva;
  reg sigmoid_table_897_0_sva;
  reg sigmoid_table_897_2_sva;
  reg sigmoid_table_125_1_sva;
  reg sigmoid_table_898_0_sva;
  reg sigmoid_table_898_2_sva;
  reg sigmoid_table_124_1_sva;
  reg sigmoid_table_899_0_sva;
  reg sigmoid_table_899_2_sva;
  reg sigmoid_table_123_1_sva;
  reg sigmoid_table_900_0_sva;
  reg sigmoid_table_900_2_sva;
  reg sigmoid_table_122_1_sva;
  reg sigmoid_table_901_0_sva;
  reg sigmoid_table_901_2_sva;
  reg sigmoid_table_121_1_sva;
  reg sigmoid_table_902_0_sva;
  reg sigmoid_table_902_2_sva;
  reg sigmoid_table_120_1_sva;
  reg sigmoid_table_903_0_sva;
  reg sigmoid_table_903_2_sva;
  reg sigmoid_table_119_1_sva;
  reg sigmoid_table_904_0_sva;
  reg sigmoid_table_904_2_sva;
  reg sigmoid_table_118_1_sva;
  reg sigmoid_table_905_0_sva;
  reg sigmoid_table_905_2_sva;
  reg sigmoid_table_117_1_sva;
  reg sigmoid_table_906_0_sva;
  reg sigmoid_table_906_2_sva;
  reg sigmoid_table_116_1_sva;
  reg sigmoid_table_907_0_sva;
  reg sigmoid_table_907_2_sva;
  reg sigmoid_table_115_1_sva;
  reg sigmoid_table_908_0_sva;
  reg sigmoid_table_908_2_sva;
  reg sigmoid_table_114_1_sva;
  reg sigmoid_table_909_0_sva;
  reg sigmoid_table_909_2_sva;
  reg sigmoid_table_113_1_sva;
  reg sigmoid_table_910_0_sva;
  reg sigmoid_table_910_2_sva;
  reg sigmoid_table_112_0_sva;
  reg sigmoid_table_911_1_sva;
  reg sigmoid_table_111_0_sva;
  reg sigmoid_table_912_1_sva;
  reg sigmoid_table_110_0_sva;
  reg sigmoid_table_913_1_sva;
  reg sigmoid_table_109_0_sva;
  reg sigmoid_table_914_1_sva;
  reg sigmoid_table_108_0_sva;
  reg sigmoid_table_915_1_sva;
  reg sigmoid_table_107_0_sva;
  reg sigmoid_table_916_1_sva;
  reg sigmoid_table_106_0_sva;
  reg sigmoid_table_917_1_sva;
  reg sigmoid_table_105_0_sva;
  reg sigmoid_table_918_1_sva;
  reg sigmoid_table_104_0_sva;
  reg sigmoid_table_919_1_sva;
  reg sigmoid_table_103_0_sva;
  reg sigmoid_table_920_1_sva;
  reg sigmoid_table_102_0_sva;
  reg sigmoid_table_921_1_sva;
  reg sigmoid_table_101_0_sva;
  reg sigmoid_table_922_1_sva;
  reg sigmoid_table_100_0_sva;
  reg sigmoid_table_923_1_sva;
  reg sigmoid_table_99_0_sva;
  reg sigmoid_table_924_1_sva;
  reg sigmoid_table_98_0_sva;
  reg sigmoid_table_925_1_sva;
  reg sigmoid_table_97_0_sva;
  reg sigmoid_table_926_1_sva;
  reg sigmoid_table_96_0_sva;
  reg sigmoid_table_927_1_sva;
  reg sigmoid_table_95_0_sva;
  reg sigmoid_table_928_1_sva;
  reg sigmoid_table_94_0_sva;
  reg sigmoid_table_929_1_sva;
  reg sigmoid_table_93_0_sva;
  reg sigmoid_table_930_1_sva;
  reg sigmoid_table_92_0_sva;
  reg sigmoid_table_931_1_sva;
  reg sigmoid_table_91_0_sva;
  reg sigmoid_table_932_1_sva;
  reg sigmoid_table_90_0_sva;
  reg sigmoid_table_933_1_sva;
  reg sigmoid_table_89_0_sva;
  reg sigmoid_table_934_1_sva;
  reg sigmoid_table_88_0_sva;
  reg sigmoid_table_935_1_sva;
  reg sigmoid_table_87_0_sva;
  reg sigmoid_table_936_1_sva;
  reg sigmoid_table_86_0_sva;
  reg sigmoid_table_937_1_sva;
  reg sigmoid_table_85_0_sva;
  reg sigmoid_table_938_1_sva;
  reg sigmoid_table_84_0_sva;
  reg sigmoid_table_939_1_sva;
  reg sigmoid_table_83_0_sva;
  reg sigmoid_table_940_1_sva;
  reg sigmoid_table_82_0_sva;
  reg sigmoid_table_941_1_sva;
  reg sigmoid_table_81_0_sva;
  reg sigmoid_table_942_1_sva;
  reg sigmoid_table_80_0_sva;
  reg sigmoid_table_943_1_sva;
  reg sigmoid_table_79_0_sva;
  reg sigmoid_table_944_1_sva;
  reg sigmoid_table_78_0_sva;
  reg sigmoid_table_945_1_sva;
  reg sigmoid_table_77_0_sva;
  reg sigmoid_table_946_1_sva;
  reg sigmoid_table_76_0_sva;
  reg sigmoid_table_947_1_sva;
  reg sigmoid_table_75_0_sva;
  reg sigmoid_table_948_1_sva;
  reg sigmoid_table_74_0_sva;
  reg sigmoid_table_949_1_sva;
  reg sigmoid_table_73_0_sva;
  reg sigmoid_table_950_1_sva;
  reg sigmoid_table_72_0_sva;
  reg sigmoid_table_951_1_sva;
  reg sigmoid_table_71_0_sva;
  reg sigmoid_table_952_1_sva;
  reg sigmoid_table_70_0_sva;
  reg sigmoid_table_953_1_sva;
  reg sigmoid_table_69_0_sva;
  reg sigmoid_table_954_1_sva;
  reg sigmoid_table_955_0_sva;
  reg sigmoid_table_956_0_sva;
  reg sigmoid_table_957_0_sva;
  reg sigmoid_table_958_0_sva;
  reg sigmoid_table_959_0_sva;
  reg sigmoid_table_960_0_sva;
  reg sigmoid_table_961_0_sva;
  reg sigmoid_table_962_0_sva;
  reg sigmoid_table_963_0_sva;
  reg sigmoid_table_964_0_sva;
  reg sigmoid_table_965_0_sva;
  reg sigmoid_table_966_0_sva;
  reg sigmoid_table_967_0_sva;
  reg sigmoid_table_968_0_sva;
  reg sigmoid_table_969_0_sva;
  reg sigmoid_table_970_0_sva;
  reg sigmoid_table_971_0_sva;
  reg sigmoid_table_972_0_sva;
  reg sigmoid_table_973_0_sva;
  reg sigmoid_table_974_0_sva;
  reg sigmoid_table_975_0_sva;
  reg sigmoid_table_976_0_sva;
  reg sigmoid_table_977_0_sva;
  reg sigmoid_table_978_0_sva;
  reg sigmoid_table_979_0_sva;
  reg sigmoid_table_980_0_sva;
  reg sigmoid_table_981_0_sva;
  reg sigmoid_table_982_0_sva;
  reg sigmoid_table_983_0_sva;
  reg sigmoid_table_984_0_sva;
  reg sigmoid_table_985_0_sva;
  reg sigmoid_table_986_0_sva;
  reg sigmoid_table_987_0_sva;
  reg sigmoid_table_988_0_sva;
  reg sigmoid_table_989_0_sva;
  reg sigmoid_table_990_0_sva;
  reg sigmoid_table_991_0_sva;
  reg sigmoid_table_992_0_sva;
  reg sigmoid_table_993_0_sva;
  reg sigmoid_table_994_0_sva;
  reg sigmoid_table_995_0_sva;
  reg sigmoid_table_996_0_sva;
  reg sigmoid_table_997_0_sva;
  reg sigmoid_table_998_0_sva;
  reg sigmoid_table_999_0_sva;
  reg sigmoid_table_1000_0_sva;
  reg sigmoid_table_1001_0_sva;
  reg sigmoid_table_1002_0_sva;
  reg sigmoid_table_1003_0_sva;
  reg sigmoid_table_1004_0_sva;
  reg sigmoid_table_1005_0_sva;
  reg sigmoid_table_1006_0_sva;
  reg sigmoid_table_1007_0_sva;
  reg sigmoid_table_1008_0_sva;
  reg sigmoid_table_1009_0_sva;
  reg sigmoid_table_1010_0_sva;
  reg sigmoid_table_1011_0_sva;
  reg sigmoid_table_1012_0_sva;
  reg sigmoid_table_1013_0_sva;
  reg sigmoid_table_1014_0_sva;
  reg sigmoid_table_1015_0_sva;
  reg sigmoid_table_1016_0_sva;
  reg sigmoid_table_1017_0_sva;
  reg sigmoid_table_1018_0_sva;
  reg sigmoid_table_1019_0_sva;
  reg sigmoid_table_1020_0_sva;
  reg sigmoid_table_1021_0_sva;
  reg sigmoid_table_1022_0_sva;
  reg sigmoid_table_1023_0_sva;
  wire sigmoid_table_69_0_sva_dfm_1;
  wire sigmoid_table_70_0_sva_dfm_1;
  wire sigmoid_table_71_0_sva_dfm_1;
  wire sigmoid_table_72_0_sva_dfm_1;
  wire sigmoid_table_73_0_sva_dfm_1;
  wire sigmoid_table_74_0_sva_dfm_1;
  wire sigmoid_table_75_0_sva_dfm_1;
  wire sigmoid_table_76_0_sva_dfm_1;
  wire sigmoid_table_77_0_sva_dfm_1;
  wire sigmoid_table_78_0_sva_dfm_1;
  wire sigmoid_table_79_0_sva_dfm_1;
  wire sigmoid_table_80_0_sva_dfm_1;
  wire sigmoid_table_81_0_sva_dfm_1;
  wire sigmoid_table_82_0_sva_dfm_1;
  wire sigmoid_table_83_0_sva_dfm_1;
  wire sigmoid_table_84_0_sva_dfm_1;
  wire sigmoid_table_85_0_sva_dfm_1;
  wire sigmoid_table_86_0_sva_dfm_1;
  wire sigmoid_table_87_0_sva_dfm_1;
  wire sigmoid_table_88_0_sva_dfm_1;
  wire sigmoid_table_89_0_sva_dfm_1;
  wire sigmoid_table_90_0_sva_dfm_1;
  wire sigmoid_table_91_0_sva_dfm_1;
  wire sigmoid_table_92_0_sva_dfm_1;
  wire sigmoid_table_93_0_sva_dfm_1;
  wire sigmoid_table_94_0_sva_dfm_1;
  wire sigmoid_table_95_0_sva_dfm_1;
  wire sigmoid_table_96_0_sva_dfm_1;
  wire sigmoid_table_97_0_sva_dfm_1;
  wire sigmoid_table_98_0_sva_dfm_1;
  wire sigmoid_table_99_0_sva_dfm_1;
  wire sigmoid_table_100_0_sva_dfm_1;
  wire sigmoid_table_101_0_sva_dfm_1;
  wire sigmoid_table_102_0_sva_dfm_1;
  wire sigmoid_table_103_0_sva_dfm_1;
  wire sigmoid_table_104_0_sva_dfm_1;
  wire sigmoid_table_105_0_sva_dfm_1;
  wire sigmoid_table_106_0_sva_dfm_1;
  wire sigmoid_table_107_0_sva_dfm_1;
  wire sigmoid_table_108_0_sva_dfm_1;
  wire sigmoid_table_109_0_sva_dfm_1;
  wire sigmoid_table_110_0_sva_dfm_1;
  wire sigmoid_table_111_0_sva_dfm_1;
  wire sigmoid_table_112_0_sva_dfm_1;
  wire sigmoid_table_139_0_sva_dfm_1;
  wire sigmoid_table_140_0_sva_dfm_1;
  wire sigmoid_table_141_0_sva_dfm_1;
  wire sigmoid_table_142_0_sva_dfm_1;
  wire sigmoid_table_143_0_sva_dfm_1;
  wire sigmoid_table_144_0_sva_dfm_1;
  wire sigmoid_table_145_0_sva_dfm_1;
  wire sigmoid_table_146_0_sva_dfm_1;
  wire sigmoid_table_147_0_sva_dfm_1;
  wire sigmoid_table_148_0_sva_dfm_1;
  wire sigmoid_table_149_0_sva_dfm_1;
  wire sigmoid_table_150_0_sva_dfm_1;
  wire sigmoid_table_151_0_sva_dfm_1;
  wire sigmoid_table_152_0_sva_dfm_1;
  wire sigmoid_table_153_0_sva_dfm_1;
  wire sigmoid_table_154_0_sva_dfm_1;
  wire sigmoid_table_155_0_sva_dfm_1;
  wire sigmoid_table_156_0_sva_dfm_1;
  wire sigmoid_table_157_0_sva_dfm_1;
  wire sigmoid_table_172_0_sva_dfm_1;
  wire sigmoid_table_173_0_sva_dfm_1;
  wire sigmoid_table_174_0_sva_dfm_1;
  wire sigmoid_table_175_0_sva_dfm_1;
  wire sigmoid_table_176_0_sva_dfm_1;
  wire sigmoid_table_177_0_sva_dfm_1;
  wire sigmoid_table_178_0_sva_dfm_1;
  wire sigmoid_table_179_0_sva_dfm_1;
  wire sigmoid_table_180_0_sva_dfm_1;
  wire sigmoid_table_181_0_sva_dfm_1;
  wire sigmoid_table_182_0_sva_dfm_1;
  wire sigmoid_table_183_0_sva_dfm_1;
  wire sigmoid_table_194_0_sva_dfm_1;
  wire sigmoid_table_195_0_sva_dfm_1;
  wire sigmoid_table_196_0_sva_dfm_1;
  wire sigmoid_table_197_0_sva_dfm_1;
  wire sigmoid_table_198_0_sva_dfm_1;
  wire sigmoid_table_199_0_sva_dfm_1;
  wire sigmoid_table_200_0_sva_dfm_1;
  wire sigmoid_table_201_0_sva_dfm_1;
  wire sigmoid_table_210_0_sva_dfm_1;
  wire sigmoid_table_211_0_sva_dfm_1;
  wire sigmoid_table_212_0_sva_dfm_1;
  wire sigmoid_table_213_0_sva_dfm_1;
  wire sigmoid_table_214_0_sva_dfm_1;
  wire sigmoid_table_215_0_sva_dfm_1;
  wire sigmoid_table_216_0_sva_dfm_1;
  wire sigmoid_table_223_0_sva_dfm_1;
  wire sigmoid_table_224_0_sva_dfm_1;
  wire sigmoid_table_225_0_sva_dfm_1;
  wire sigmoid_table_226_0_sva_dfm_1;
  wire sigmoid_table_227_0_sva_dfm_1;
  wire sigmoid_table_228_0_sva_dfm_1;
  wire sigmoid_table_234_0_sva_dfm_1;
  wire sigmoid_table_235_0_sva_dfm_1;
  wire sigmoid_table_236_0_sva_dfm_1;
  wire sigmoid_table_237_0_sva_dfm_1;
  wire sigmoid_table_238_0_sva_dfm_1;
  wire sigmoid_table_243_0_sva_dfm_1;
  wire sigmoid_table_244_0_sva_dfm_1;
  wire sigmoid_table_245_0_sva_dfm_1;
  wire sigmoid_table_246_0_sva_dfm_1;
  wire sigmoid_table_251_0_sva_dfm_1;
  wire sigmoid_table_252_0_sva_dfm_1;
  wire sigmoid_table_253_0_sva_dfm_1;
  wire sigmoid_table_254_0_sva_dfm_1;
  wire sigmoid_table_259_0_sva_dfm_1;
  wire sigmoid_table_260_0_sva_dfm_1;
  wire sigmoid_table_261_0_sva_dfm_1;
  wire sigmoid_table_265_0_sva_dfm_1;
  wire sigmoid_table_266_0_sva_dfm_1;
  wire sigmoid_table_267_0_sva_dfm_1;
  wire sigmoid_table_271_0_sva_dfm_1;
  wire sigmoid_table_272_0_sva_dfm_1;
  wire sigmoid_table_273_0_sva_dfm_1;
  wire sigmoid_table_276_0_sva_dfm_1;
  wire sigmoid_table_277_0_sva_dfm_1;
  wire sigmoid_table_278_0_sva_dfm_1;
  wire sigmoid_table_282_0_sva_dfm_1;
  wire sigmoid_table_283_0_sva_dfm_1;
  wire sigmoid_table_286_0_sva_dfm_1;
  wire sigmoid_table_287_0_sva_dfm_1;
  wire sigmoid_table_291_0_sva_dfm_1;
  wire sigmoid_table_292_0_sva_dfm_1;
  wire sigmoid_table_295_0_sva_dfm_1;
  wire sigmoid_table_296_0_sva_dfm_1;
  wire sigmoid_table_299_0_sva_dfm_1;
  wire sigmoid_table_300_0_sva_dfm_1;
  wire sigmoid_table_302_0_sva_dfm_1;
  wire sigmoid_table_303_0_sva_dfm_1;
  wire sigmoid_table_306_0_sva_dfm_1;
  wire sigmoid_table_307_0_sva_dfm_1;
  wire sigmoid_table_309_0_sva_dfm_1;
  wire sigmoid_table_310_0_sva_dfm_1;
  wire sigmoid_table_312_0_sva_dfm_1;
  wire sigmoid_table_313_0_sva_dfm_1;
  wire sigmoid_table_315_0_sva_dfm_1;
  wire sigmoid_table_316_0_sva_dfm_1;
  wire sigmoid_table_318_0_sva_dfm_1;
  wire sigmoid_table_319_0_sva_dfm_1;
  wire sigmoid_table_321_0_sva_dfm_1;
  wire sigmoid_table_324_0_sva_dfm_1;
  wire sigmoid_table_326_0_sva_dfm_1;
  wire sigmoid_table_327_0_sva_dfm_1;
  wire sigmoid_table_329_0_sva_dfm_1;
  wire sigmoid_table_331_0_sva_dfm_1;
  wire sigmoid_table_334_0_sva_dfm_1;
  wire sigmoid_table_336_0_sva_dfm_1;
  wire sigmoid_table_338_0_sva_dfm_1;
  wire sigmoid_table_340_0_sva_dfm_1;
  wire sigmoid_table_342_0_sva_dfm_1;
  wire sigmoid_table_344_0_sva_dfm_1;
  wire sigmoid_table_346_0_sva_dfm_1;
  wire sigmoid_table_348_0_sva_dfm_1;
  wire sigmoid_table_350_0_sva_dfm_1;
  wire sigmoid_table_352_0_sva_dfm_1;
  wire sigmoid_table_354_0_sva_dfm_1;
  wire sigmoid_table_355_0_sva_dfm_1;
  wire sigmoid_table_357_0_sva_dfm_1;
  wire sigmoid_table_359_0_sva_dfm_1;
  wire sigmoid_table_360_0_sva_dfm_1;
  wire sigmoid_table_362_0_sva_dfm_1;
  wire sigmoid_table_365_0_sva_dfm_1;
  wire sigmoid_table_368_0_sva_dfm_1;
  wire sigmoid_table_369_0_sva_dfm_1;
  wire sigmoid_table_371_0_sva_dfm_1;
  wire sigmoid_table_372_0_sva_dfm_1;
  wire sigmoid_table_375_0_sva_dfm_1;
  wire sigmoid_table_376_0_sva_dfm_1;
  wire sigmoid_table_379_0_sva_dfm_1;
  wire sigmoid_table_380_0_sva_dfm_1;
  wire sigmoid_table_381_0_sva_dfm_1;
  wire sigmoid_table_385_0_sva_dfm_1;
  wire sigmoid_table_386_0_sva_dfm_1;
  wire sigmoid_table_387_0_sva_dfm_1;
  wire sigmoid_table_394_0_sva_dfm_1;
  wire sigmoid_table_395_0_sva_dfm_1;
  wire sigmoid_table_396_0_sva_dfm_1;
  wire sigmoid_table_397_0_sva_dfm_1;
  wire sigmoid_table_398_0_sva_dfm_1;
  wire sigmoid_table_399_0_sva_dfm_1;
  wire sigmoid_table_400_0_sva_dfm_1;
  wire sigmoid_table_401_0_sva_dfm_1;
  wire sigmoid_table_402_0_sva_dfm_1;
  wire sigmoid_table_403_0_sva_dfm_1;
  wire sigmoid_table_404_0_sva_dfm_1;
  wire sigmoid_table_405_0_sva_dfm_1;
  wire sigmoid_table_411_0_sva_dfm_1;
  wire sigmoid_table_412_0_sva_dfm_1;
  wire sigmoid_table_413_0_sva_dfm_1;
  wire sigmoid_table_417_0_sva_dfm_1;
  wire sigmoid_table_418_0_sva_dfm_1;
  wire sigmoid_table_421_0_sva_dfm_1;
  wire sigmoid_table_422_0_sva_dfm_1;
  wire sigmoid_table_425_0_sva_dfm_1;
  wire sigmoid_table_426_0_sva_dfm_1;
  wire sigmoid_table_428_0_sva_dfm_1;
  wire sigmoid_table_429_0_sva_dfm_1;
  wire sigmoid_table_431_0_sva_dfm_1;
  wire sigmoid_table_434_0_sva_dfm_1;
  wire sigmoid_table_436_0_sva_dfm_1;
  wire sigmoid_table_438_0_sva_dfm_1;
  wire sigmoid_table_441_0_sva_dfm_1;
  wire sigmoid_table_443_0_sva_dfm_1;
  wire sigmoid_table_446_0_sva_dfm_1;
  wire sigmoid_table_448_0_sva_dfm_1;
  wire sigmoid_table_450_0_sva_dfm_1;
  wire sigmoid_table_453_0_sva_dfm_1;
  wire sigmoid_table_455_0_sva_dfm_1;
  wire sigmoid_table_456_0_sva_dfm_1;
  wire sigmoid_table_458_0_sva_dfm_1;
  wire sigmoid_table_459_0_sva_dfm_1;
  wire sigmoid_table_462_0_sva_dfm_1;
  wire sigmoid_table_463_0_sva_dfm_1;
  wire sigmoid_table_466_0_sva_dfm_1;
  wire sigmoid_table_467_0_sva_dfm_1;
  wire sigmoid_table_470_0_sva_dfm_1;
  wire sigmoid_table_471_0_sva_dfm_1;
  wire sigmoid_table_472_0_sva_dfm_1;
  wire sigmoid_table_475_0_sva_dfm_1;
  wire sigmoid_table_476_0_sva_dfm_1;
  wire sigmoid_table_477_0_sva_dfm_1;
  wire sigmoid_table_478_0_sva_dfm_1;
  wire sigmoid_table_483_0_sva_dfm_1;
  wire sigmoid_table_484_0_sva_dfm_1;
  wire sigmoid_table_485_0_sva_dfm_1;
  wire sigmoid_table_486_0_sva_dfm_1;
  wire sigmoid_table_487_0_sva_dfm_1;
  wire sigmoid_table_488_0_sva_dfm_1;
  wire sigmoid_table_516_0_sva_dfm_1;
  wire sigmoid_table_517_0_sva_dfm_1;
  wire sigmoid_table_518_0_sva_dfm_1;
  wire sigmoid_table_519_0_sva_dfm_1;
  wire sigmoid_table_520_0_sva_dfm_1;
  wire sigmoid_table_521_0_sva_dfm_1;
  wire sigmoid_table_522_0_sva_dfm_1;
  wire sigmoid_table_523_0_sva_dfm_1;
  wire sigmoid_table_524_0_sva_dfm_1;
  wire sigmoid_table_525_0_sva_dfm_1;
  wire sigmoid_table_526_0_sva_dfm_1;
  wire sigmoid_table_527_0_sva_dfm_1;
  wire sigmoid_table_528_0_sva_dfm_1;
  wire sigmoid_table_529_0_sva_dfm_1;
  wire sigmoid_table_530_0_sva_dfm_1;
  wire sigmoid_table_531_0_sva_dfm_1;
  wire sigmoid_table_532_0_sva_dfm_1;
  wire sigmoid_table_533_0_sva_dfm_1;
  wire sigmoid_table_534_0_sva_dfm_1;
  wire sigmoid_table_535_0_sva_dfm_1;
  wire sigmoid_table_542_0_sva_dfm_1;
  wire sigmoid_table_543_0_sva_dfm_1;
  wire sigmoid_table_544_0_sva_dfm_1;
  wire sigmoid_table_545_0_sva_dfm_1;
  wire sigmoid_table_550_0_sva_dfm_1;
  wire sigmoid_table_551_0_sva_dfm_1;
  wire sigmoid_table_555_0_sva_dfm_1;
  wire sigmoid_table_556_0_sva_dfm_1;
  wire sigmoid_table_559_0_sva_dfm_1;
  wire sigmoid_table_560_0_sva_dfm_1;
  wire sigmoid_table_563_0_sva_dfm_1;
  wire sigmoid_table_564_0_sva_dfm_1;
  wire sigmoid_table_567_0_sva_dfm_1;
  wire sigmoid_table_570_0_sva_dfm_1;
  wire sigmoid_table_572_0_sva_dfm_1;
  wire sigmoid_table_573_0_sva_dfm_1;
  wire sigmoid_table_575_0_sva_dfm_1;
  wire sigmoid_table_577_0_sva_dfm_1;
  wire sigmoid_table_579_0_sva_dfm_1;
  wire sigmoid_table_580_0_sva_dfm_1;
  wire sigmoid_table_582_0_sva_dfm_1;
  wire sigmoid_table_584_0_sva_dfm_1;
  wire sigmoid_table_585_0_sva_dfm_1;
  wire sigmoid_table_587_0_sva_dfm_1;
  wire sigmoid_table_589_0_sva_dfm_1;
  wire sigmoid_table_591_0_sva_dfm_1;
  wire sigmoid_table_592_0_sva_dfm_1;
  wire sigmoid_table_594_0_sva_dfm_1;
  wire sigmoid_table_597_0_sva_dfm_1;
  wire sigmoid_table_600_0_sva_dfm_1;
  wire sigmoid_table_601_0_sva_dfm_1;
  wire sigmoid_table_604_0_sva_dfm_1;
  wire sigmoid_table_605_0_sva_dfm_1;
  wire sigmoid_table_608_0_sva_dfm_1;
  wire sigmoid_table_609_0_sva_dfm_1;
  wire sigmoid_table_610_0_sva_dfm_1;
  wire sigmoid_table_614_0_sva_dfm_1;
  wire sigmoid_table_615_0_sva_dfm_1;
  wire sigmoid_table_616_0_sva_dfm_1;
  wire sigmoid_table_617_0_sva_dfm_1;
  wire sigmoid_table_618_0_sva_dfm_1;
  wire sigmoid_table_631_0_sva_dfm_1;
  wire sigmoid_table_632_0_sva_dfm_1;
  wire sigmoid_table_633_0_sva_dfm_1;
  wire sigmoid_table_634_0_sva_dfm_1;
  wire sigmoid_table_635_0_sva_dfm_1;
  wire sigmoid_table_636_0_sva_dfm_1;
  wire sigmoid_table_640_0_sva_dfm_1;
  wire sigmoid_table_641_0_sva_dfm_1;
  wire sigmoid_table_642_0_sva_dfm_1;
  wire sigmoid_table_646_0_sva_dfm_1;
  wire sigmoid_table_647_0_sva_dfm_1;
  wire sigmoid_table_650_0_sva_dfm_1;
  wire sigmoid_table_651_0_sva_dfm_1;
  wire sigmoid_table_654_0_sva_dfm_1;
  wire sigmoid_table_657_0_sva_dfm_1;
  wire sigmoid_table_658_0_sva_dfm_1;
  wire sigmoid_table_660_0_sva_dfm_1;
  wire sigmoid_table_661_0_sva_dfm_1;
  wire sigmoid_table_663_0_sva_dfm_1;
  wire sigmoid_table_666_0_sva_dfm_1;
  wire sigmoid_table_668_0_sva_dfm_1;
  wire sigmoid_table_671_0_sva_dfm_1;
  wire sigmoid_table_673_0_sva_dfm_1;
  wire sigmoid_table_675_0_sva_dfm_1;
  wire sigmoid_table_677_0_sva_dfm_1;
  wire sigmoid_table_679_0_sva_dfm_1;
  wire sigmoid_table_681_0_sva_dfm_1;
  wire sigmoid_table_683_0_sva_dfm_1;
  wire sigmoid_table_685_0_sva_dfm_1;
  wire sigmoid_table_687_0_sva_dfm_1;
  wire sigmoid_table_689_0_sva_dfm_1;
  wire sigmoid_table_691_0_sva_dfm_1;
  wire sigmoid_table_692_0_sva_dfm_1;
  wire sigmoid_table_694_0_sva_dfm_1;
  wire sigmoid_table_696_0_sva_dfm_1;
  wire sigmoid_table_699_0_sva_dfm_1;
  wire sigmoid_table_701_0_sva_dfm_1;
  wire sigmoid_table_702_0_sva_dfm_1;
  wire sigmoid_table_704_0_sva_dfm_1;
  wire sigmoid_table_707_0_sva_dfm_1;
  wire sigmoid_table_710_0_sva_dfm_1;
  wire sigmoid_table_713_0_sva_dfm_1;
  wire sigmoid_table_716_0_sva_dfm_1;
  wire sigmoid_table_719_0_sva_dfm_1;
  wire sigmoid_table_720_0_sva_dfm_1;
  wire sigmoid_table_723_0_sva_dfm_1;
  wire sigmoid_table_726_0_sva_dfm_1;
  wire sigmoid_table_727_0_sva_dfm_1;
  wire sigmoid_table_730_0_sva_dfm_1;
  wire sigmoid_table_731_0_sva_dfm_1;
  wire sigmoid_table_734_0_sva_dfm_1;
  wire sigmoid_table_735_0_sva_dfm_1;
  wire sigmoid_table_736_0_sva_dfm_1;
  wire sigmoid_table_739_0_sva_dfm_1;
  wire sigmoid_table_740_0_sva_dfm_1;
  wire sigmoid_table_743_0_sva_dfm_1;
  wire sigmoid_table_744_0_sva_dfm_1;
  wire sigmoid_table_745_0_sva_dfm_1;
  wire sigmoid_table_748_0_sva_dfm_1;
  wire sigmoid_table_749_0_sva_dfm_1;
  wire sigmoid_table_750_0_sva_dfm_1;
  wire sigmoid_table_754_0_sva_dfm_1;
  wire sigmoid_table_755_0_sva_dfm_1;
  wire sigmoid_table_756_0_sva_dfm_1;
  wire sigmoid_table_760_0_sva_dfm_1;
  wire sigmoid_table_761_0_sva_dfm_1;
  wire sigmoid_table_762_0_sva_dfm_1;
  wire sigmoid_table_766_0_sva_dfm_1;
  wire sigmoid_table_767_0_sva_dfm_1;
  wire sigmoid_table_768_0_sva_dfm_1;
  wire sigmoid_table_769_0_sva_dfm_1;
  wire sigmoid_table_774_0_sva_dfm_1;
  wire sigmoid_table_775_0_sva_dfm_1;
  wire sigmoid_table_776_0_sva_dfm_1;
  wire sigmoid_table_777_0_sva_dfm_1;
  wire sigmoid_table_782_0_sva_dfm_1;
  wire sigmoid_table_783_0_sva_dfm_1;
  wire sigmoid_table_784_0_sva_dfm_1;
  wire sigmoid_table_785_0_sva_dfm_1;
  wire sigmoid_table_791_0_sva_dfm_1;
  wire sigmoid_table_792_0_sva_dfm_1;
  wire sigmoid_table_793_0_sva_dfm_1;
  wire sigmoid_table_794_0_sva_dfm_1;
  wire sigmoid_table_795_0_sva_dfm_1;
  wire sigmoid_table_802_0_sva_dfm_1;
  wire sigmoid_table_803_0_sva_dfm_1;
  wire sigmoid_table_804_0_sva_dfm_1;
  wire sigmoid_table_805_0_sva_dfm_1;
  wire sigmoid_table_806_0_sva_dfm_1;
  wire sigmoid_table_807_0_sva_dfm_1;
  wire sigmoid_table_815_0_sva_dfm_1;
  wire sigmoid_table_816_0_sva_dfm_1;
  wire sigmoid_table_817_0_sva_dfm_1;
  wire sigmoid_table_818_0_sva_dfm_1;
  wire sigmoid_table_819_0_sva_dfm_1;
  wire sigmoid_table_820_0_sva_dfm_1;
  wire sigmoid_table_821_0_sva_dfm_1;
  wire sigmoid_table_831_0_sva_dfm_1;
  wire sigmoid_table_832_0_sva_dfm_1;
  wire sigmoid_table_833_0_sva_dfm_1;
  wire sigmoid_table_834_0_sva_dfm_1;
  wire sigmoid_table_835_0_sva_dfm_1;
  wire sigmoid_table_836_0_sva_dfm_1;
  wire sigmoid_table_837_0_sva_dfm_1;
  wire sigmoid_table_838_0_sva_dfm_1;
  wire sigmoid_table_839_0_sva_dfm_1;
  wire sigmoid_table_840_0_sva_dfm_1;
  wire sigmoid_table_853_0_sva_dfm_1;
  wire sigmoid_table_854_0_sva_dfm_1;
  wire sigmoid_table_855_0_sva_dfm_1;
  wire sigmoid_table_856_0_sva_dfm_1;
  wire sigmoid_table_857_0_sva_dfm_1;
  wire sigmoid_table_858_0_sva_dfm_1;
  wire sigmoid_table_859_0_sva_dfm_1;
  wire sigmoid_table_860_0_sva_dfm_1;
  wire sigmoid_table_861_0_sva_dfm_1;
  wire sigmoid_table_862_0_sva_dfm_1;
  wire sigmoid_table_863_0_sva_dfm_1;
  wire sigmoid_table_864_0_sva_dfm_1;
  wire sigmoid_table_865_0_sva_dfm_1;
  wire sigmoid_table_866_0_sva_dfm_1;
  wire sigmoid_table_885_0_sva_dfm_1;
  wire sigmoid_table_886_0_sva_dfm_1;
  wire sigmoid_table_887_0_sva_dfm_1;
  wire sigmoid_table_888_0_sva_dfm_1;
  wire sigmoid_table_889_0_sva_dfm_1;
  wire sigmoid_table_890_0_sva_dfm_1;
  wire sigmoid_table_891_0_sva_dfm_1;
  wire sigmoid_table_892_0_sva_dfm_1;
  wire sigmoid_table_893_0_sva_dfm_1;
  wire sigmoid_table_894_0_sva_dfm_1;
  wire sigmoid_table_895_0_sva_dfm_1;
  wire sigmoid_table_896_0_sva_dfm_1;
  wire sigmoid_table_897_0_sva_dfm_1;
  wire sigmoid_table_898_0_sva_dfm_1;
  wire sigmoid_table_899_0_sva_dfm_1;
  wire sigmoid_table_900_0_sva_dfm_1;
  wire sigmoid_table_901_0_sva_dfm_1;
  wire sigmoid_table_902_0_sva_dfm_1;
  wire sigmoid_table_903_0_sva_dfm_1;
  wire sigmoid_table_904_0_sva_dfm_1;
  wire sigmoid_table_905_0_sva_dfm_1;
  wire sigmoid_table_906_0_sva_dfm_1;
  wire sigmoid_table_907_0_sva_dfm_1;
  wire sigmoid_table_908_0_sva_dfm_1;
  wire sigmoid_table_909_0_sva_dfm_1;
  wire sigmoid_table_910_0_sva_dfm_1;
  wire sigmoid_table_955_0_sva_dfm_1;
  wire sigmoid_table_956_0_sva_dfm_1;
  wire sigmoid_table_957_0_sva_dfm_1;
  wire sigmoid_table_958_0_sva_dfm_1;
  wire sigmoid_table_959_0_sva_dfm_1;
  wire sigmoid_table_960_0_sva_dfm_1;
  wire sigmoid_table_961_0_sva_dfm_1;
  wire sigmoid_table_962_0_sva_dfm_1;
  wire sigmoid_table_963_0_sva_dfm_1;
  wire sigmoid_table_964_0_sva_dfm_1;
  wire sigmoid_table_965_0_sva_dfm_1;
  wire sigmoid_table_966_0_sva_dfm_1;
  wire sigmoid_table_967_0_sva_dfm_1;
  wire sigmoid_table_968_0_sva_dfm_1;
  wire sigmoid_table_969_0_sva_dfm_1;
  wire sigmoid_table_970_0_sva_dfm_1;
  wire sigmoid_table_971_0_sva_dfm_1;
  wire sigmoid_table_972_0_sva_dfm_1;
  wire sigmoid_table_973_0_sva_dfm_1;
  wire sigmoid_table_974_0_sva_dfm_1;
  wire sigmoid_table_975_0_sva_dfm_1;
  wire sigmoid_table_976_0_sva_dfm_1;
  wire sigmoid_table_977_0_sva_dfm_1;
  wire sigmoid_table_978_0_sva_dfm_1;
  wire sigmoid_table_979_0_sva_dfm_1;
  wire sigmoid_table_980_0_sva_dfm_1;
  wire sigmoid_table_981_0_sva_dfm_1;
  wire sigmoid_table_982_0_sva_dfm_1;
  wire sigmoid_table_983_0_sva_dfm_1;
  wire sigmoid_table_984_0_sva_dfm_1;
  wire sigmoid_table_985_0_sva_dfm_1;
  wire sigmoid_table_986_0_sva_dfm_1;
  wire sigmoid_table_987_0_sva_dfm_1;
  wire sigmoid_table_988_0_sva_dfm_1;
  wire sigmoid_table_989_0_sva_dfm_1;
  wire sigmoid_table_990_0_sva_dfm_1;
  wire sigmoid_table_991_0_sva_dfm_1;
  wire sigmoid_table_992_0_sva_dfm_1;
  wire sigmoid_table_993_0_sva_dfm_1;
  wire sigmoid_table_994_0_sva_dfm_1;
  wire sigmoid_table_995_0_sva_dfm_1;
  wire sigmoid_table_996_0_sva_dfm_1;
  wire sigmoid_table_997_0_sva_dfm_1;
  wire sigmoid_table_998_0_sva_dfm_1;
  wire sigmoid_table_999_0_sva_dfm_1;
  wire sigmoid_table_1000_0_sva_dfm_1;
  wire sigmoid_table_1001_0_sva_dfm_1;
  wire sigmoid_table_1002_0_sva_dfm_1;
  wire sigmoid_table_1003_0_sva_dfm_1;
  wire sigmoid_table_1004_0_sva_dfm_1;
  wire sigmoid_table_1005_0_sva_dfm_1;
  wire sigmoid_table_1006_0_sva_dfm_1;
  wire sigmoid_table_1007_0_sva_dfm_1;
  wire sigmoid_table_1008_0_sva_dfm_1;
  wire sigmoid_table_1009_0_sva_dfm_1;
  wire sigmoid_table_1010_0_sva_dfm_1;
  wire sigmoid_table_1011_0_sva_dfm_1;
  wire sigmoid_table_1012_0_sva_dfm_1;
  wire sigmoid_table_1013_0_sva_dfm_1;
  wire sigmoid_table_1014_0_sva_dfm_1;
  wire sigmoid_table_1015_0_sva_dfm_1;
  wire sigmoid_table_1016_0_sva_dfm_1;
  wire sigmoid_table_1017_0_sva_dfm_1;
  wire sigmoid_table_1018_0_sva_dfm_1;
  wire sigmoid_table_1019_0_sva_dfm_1;
  wire sigmoid_table_1020_0_sva_dfm_1;
  wire sigmoid_table_1021_0_sva_dfm_1;
  wire sigmoid_table_1022_0_sva_dfm_1;
  wire sigmoid_table_1023_0_sva_dfm_1;
  wire sigmoid_table_512_9_sva_dfm_1;
  wire sigmoid_table_513_9_sva_dfm_1;
  wire sigmoid_table_514_9_sva_dfm_1;
  wire sigmoid_table_515_9_sva_dfm_1;
  wire sigmoid_table_516_9_sva_dfm_1;
  wire sigmoid_table_517_9_sva_dfm_1;
  wire sigmoid_table_518_9_sva_dfm_1;
  wire sigmoid_table_519_9_sva_dfm_1;
  wire sigmoid_table_520_9_sva_dfm_1;
  wire sigmoid_table_521_9_sva_dfm_1;
  wire sigmoid_table_522_9_sva_dfm_1;
  wire sigmoid_table_523_9_sva_dfm_1;
  wire sigmoid_table_524_9_sva_dfm_1;
  wire sigmoid_table_525_9_sva_dfm_1;
  wire sigmoid_table_526_9_sva_dfm_1;
  wire sigmoid_table_527_9_sva_dfm_1;
  wire sigmoid_table_528_9_sva_dfm_1;
  wire sigmoid_table_529_9_sva_dfm_1;
  wire sigmoid_table_530_9_sva_dfm_1;
  wire sigmoid_table_531_9_sva_dfm_1;
  wire sigmoid_table_532_9_sva_dfm_1;
  wire sigmoid_table_533_9_sva_dfm_1;
  wire sigmoid_table_534_9_sva_dfm_1;
  wire sigmoid_table_535_9_sva_dfm_1;
  wire sigmoid_table_536_9_sva_dfm_1;
  wire sigmoid_table_537_9_sva_dfm_1;
  wire sigmoid_table_538_9_sva_dfm_1;
  wire sigmoid_table_539_9_sva_dfm_1;
  wire sigmoid_table_540_9_sva_dfm_1;
  wire sigmoid_table_541_9_sva_dfm_1;
  wire sigmoid_table_542_9_sva_dfm_1;
  wire sigmoid_table_543_9_sva_dfm_1;
  wire sigmoid_table_544_9_sva_dfm_1;
  wire sigmoid_table_545_9_sva_dfm_1;
  wire sigmoid_table_546_9_sva_dfm_1;
  wire sigmoid_table_547_9_sva_dfm_1;
  wire sigmoid_table_548_9_sva_dfm_1;
  wire sigmoid_table_549_9_sva_dfm_1;
  wire sigmoid_table_550_9_sva_dfm_1;
  wire sigmoid_table_551_9_sva_dfm_1;
  wire sigmoid_table_552_9_sva_dfm_1;
  wire sigmoid_table_553_9_sva_dfm_1;
  wire sigmoid_table_554_9_sva_dfm_1;
  wire sigmoid_table_555_9_sva_dfm_1;
  wire sigmoid_table_556_9_sva_dfm_1;
  wire sigmoid_table_557_9_sva_dfm_1;
  wire sigmoid_table_558_9_sva_dfm_1;
  wire sigmoid_table_559_9_sva_dfm_1;
  wire sigmoid_table_560_9_sva_dfm_1;
  wire sigmoid_table_561_9_sva_dfm_1;
  wire sigmoid_table_562_9_sva_dfm_1;
  wire sigmoid_table_563_9_sva_dfm_1;
  wire sigmoid_table_564_9_sva_dfm_1;
  wire sigmoid_table_565_9_sva_dfm_1;
  wire sigmoid_table_566_9_sva_dfm_1;
  wire sigmoid_table_567_9_sva_dfm_1;
  wire sigmoid_table_568_9_sva_dfm_1;
  wire sigmoid_table_569_9_sva_dfm_1;
  wire sigmoid_table_570_9_sva_dfm_1;
  wire sigmoid_table_571_9_sva_dfm_1;
  wire sigmoid_table_572_9_sva_dfm_1;
  wire sigmoid_table_573_9_sva_dfm_1;
  wire sigmoid_table_574_9_sva_dfm_1;
  wire sigmoid_table_575_9_sva_dfm_1;
  wire sigmoid_table_576_9_sva_dfm_1;
  wire sigmoid_table_577_9_sva_dfm_1;
  wire sigmoid_table_578_9_sva_dfm_1;
  wire sigmoid_table_579_9_sva_dfm_1;
  wire sigmoid_table_580_9_sva_dfm_1;
  wire sigmoid_table_581_9_sva_dfm_1;
  wire sigmoid_table_582_9_sva_dfm_1;
  wire sigmoid_table_583_8_sva_dfm_1;
  wire sigmoid_table_584_8_sva_dfm_1;
  wire sigmoid_table_585_8_sva_dfm_1;
  wire sigmoid_table_586_8_sva_dfm_1;
  wire sigmoid_table_587_8_sva_dfm_1;
  wire sigmoid_table_588_8_sva_dfm_1;
  wire sigmoid_table_589_8_sva_dfm_1;
  wire sigmoid_table_590_8_sva_dfm_1;
  wire sigmoid_table_591_8_sva_dfm_1;
  wire sigmoid_table_592_8_sva_dfm_1;
  wire sigmoid_table_593_8_sva_dfm_1;
  wire sigmoid_table_594_8_sva_dfm_1;
  wire sigmoid_table_595_8_sva_dfm_1;
  wire sigmoid_table_596_8_sva_dfm_1;
  wire sigmoid_table_597_8_sva_dfm_1;
  wire sigmoid_table_598_8_sva_dfm_1;
  wire sigmoid_table_599_8_sva_dfm_1;
  wire sigmoid_table_600_8_sva_dfm_1;
  wire sigmoid_table_601_8_sva_dfm_1;
  wire sigmoid_table_602_8_sva_dfm_1;
  wire sigmoid_table_603_8_sva_dfm_1;
  wire sigmoid_table_604_8_sva_dfm_1;
  wire sigmoid_table_605_8_sva_dfm_1;
  wire sigmoid_table_606_8_sva_dfm_1;
  wire sigmoid_table_607_8_sva_dfm_1;
  wire sigmoid_table_608_8_sva_dfm_1;
  wire sigmoid_table_609_8_sva_dfm_1;
  wire sigmoid_table_610_8_sva_dfm_1;
  wire sigmoid_table_611_8_sva_dfm_1;
  wire sigmoid_table_612_8_sva_dfm_1;
  wire sigmoid_table_613_8_sva_dfm_1;
  wire sigmoid_table_614_8_sva_dfm_1;
  wire sigmoid_table_615_8_sva_dfm_1;
  wire sigmoid_table_616_8_sva_dfm_1;
  wire sigmoid_table_617_8_sva_dfm_1;
  wire sigmoid_table_618_8_sva_dfm_1;
  wire sigmoid_table_619_8_sva_dfm_1;
  wire sigmoid_table_620_8_sva_dfm_1;
  wire sigmoid_table_621_8_sva_dfm_1;
  wire sigmoid_table_622_8_sva_dfm_1;
  wire sigmoid_table_623_8_sva_dfm_1;
  wire sigmoid_table_624_8_sva_dfm_1;
  wire sigmoid_table_625_8_sva_dfm_1;
  wire sigmoid_table_626_8_sva_dfm_1;
  wire sigmoid_table_627_8_sva_dfm_1;
  wire sigmoid_table_628_8_sva_dfm_1;
  wire sigmoid_table_629_8_sva_dfm_1;
  wire sigmoid_table_630_8_sva_dfm_1;
  wire sigmoid_table_631_8_sva_dfm_1;
  wire sigmoid_table_632_8_sva_dfm_1;
  wire sigmoid_table_633_8_sva_dfm_1;
  wire sigmoid_table_634_8_sva_dfm_1;
  wire sigmoid_table_635_8_sva_dfm_1;
  wire sigmoid_table_636_8_sva_dfm_1;
  wire sigmoid_table_637_7_sva_dfm_1;
  wire sigmoid_table_638_7_sva_dfm_1;
  wire sigmoid_table_639_7_sva_dfm_1;
  wire sigmoid_table_640_7_sva_dfm_1;
  wire sigmoid_table_641_7_sva_dfm_1;
  wire sigmoid_table_642_7_sva_dfm_1;
  wire sigmoid_table_643_7_sva_dfm_1;
  wire sigmoid_table_644_7_sva_dfm_1;
  wire sigmoid_table_645_7_sva_dfm_1;
  wire sigmoid_table_646_7_sva_dfm_1;
  wire sigmoid_table_647_7_sva_dfm_1;
  wire sigmoid_table_648_7_sva_dfm_1;
  wire sigmoid_table_649_7_sva_dfm_1;
  wire sigmoid_table_650_7_sva_dfm_1;
  wire sigmoid_table_651_7_sva_dfm_1;
  wire sigmoid_table_652_7_sva_dfm_1;
  wire sigmoid_table_653_7_sva_dfm_1;
  wire sigmoid_table_654_7_sva_dfm_1;
  wire sigmoid_table_655_7_sva_dfm_1;
  wire sigmoid_table_656_7_sva_dfm_1;
  wire sigmoid_table_657_7_sva_dfm_1;
  wire sigmoid_table_658_7_sva_dfm_1;
  wire sigmoid_table_659_7_sva_dfm_1;
  wire sigmoid_table_660_7_sva_dfm_1;
  wire sigmoid_table_661_7_sva_dfm_1;
  wire sigmoid_table_662_7_sva_dfm_1;
  wire sigmoid_table_663_7_sva_dfm_1;
  wire sigmoid_table_664_7_sva_dfm_1;
  wire sigmoid_table_665_7_sva_dfm_1;
  wire sigmoid_table_666_7_sva_dfm_1;
  wire sigmoid_table_667_7_sva_dfm_1;
  wire sigmoid_table_668_7_sva_dfm_1;
  wire sigmoid_table_669_7_sva_dfm_1;
  wire sigmoid_table_670_7_sva_dfm_1;
  wire sigmoid_table_671_7_sva_dfm_1;
  wire sigmoid_table_672_7_sva_dfm_1;
  wire sigmoid_table_673_7_sva_dfm_1;
  wire sigmoid_table_674_7_sva_dfm_1;
  wire sigmoid_table_675_7_sva_dfm_1;
  wire sigmoid_table_676_7_sva_dfm_1;
  wire sigmoid_table_677_7_sva_dfm_1;
  wire sigmoid_table_678_7_sva_dfm_1;
  wire sigmoid_table_679_7_sva_dfm_1;
  wire sigmoid_table_680_7_sva_dfm_1;
  wire sigmoid_table_681_7_sva_dfm_1;
  wire sigmoid_table_682_7_sva_dfm_1;
  wire sigmoid_table_683_7_sva_dfm_1;
  wire sigmoid_table_684_7_sva_dfm_1;
  wire sigmoid_table_685_7_sva_dfm_1;
  wire sigmoid_table_686_6_sva_dfm_1;
  wire sigmoid_table_687_6_sva_dfm_1;
  wire sigmoid_table_688_6_sva_dfm_1;
  wire sigmoid_table_689_6_sva_dfm_1;
  wire sigmoid_table_690_6_sva_dfm_1;
  wire sigmoid_table_691_6_sva_dfm_1;
  wire sigmoid_table_692_6_sva_dfm_1;
  wire sigmoid_table_693_6_sva_dfm_1;
  wire sigmoid_table_694_6_sva_dfm_1;
  wire sigmoid_table_695_6_sva_dfm_1;
  wire sigmoid_table_696_6_sva_dfm_1;
  wire sigmoid_table_697_6_sva_dfm_1;
  wire sigmoid_table_698_6_sva_dfm_1;
  wire sigmoid_table_699_6_sva_dfm_1;
  wire sigmoid_table_700_6_sva_dfm_1;
  wire sigmoid_table_701_6_sva_dfm_1;
  wire sigmoid_table_702_6_sva_dfm_1;
  wire sigmoid_table_703_6_sva_dfm_1;
  wire sigmoid_table_704_6_sva_dfm_1;
  wire sigmoid_table_705_6_sva_dfm_1;
  wire sigmoid_table_706_6_sva_dfm_1;
  wire sigmoid_table_707_6_sva_dfm_1;
  wire sigmoid_table_708_6_sva_dfm_1;
  wire sigmoid_table_709_6_sva_dfm_1;
  wire sigmoid_table_710_6_sva_dfm_1;
  wire sigmoid_table_711_6_sva_dfm_1;
  wire sigmoid_table_712_6_sva_dfm_1;
  wire sigmoid_table_713_6_sva_dfm_1;
  wire sigmoid_table_714_6_sva_dfm_1;
  wire sigmoid_table_715_6_sva_dfm_1;
  wire sigmoid_table_716_6_sva_dfm_1;
  wire sigmoid_table_717_6_sva_dfm_1;
  wire sigmoid_table_718_6_sva_dfm_1;
  wire sigmoid_table_719_6_sva_dfm_1;
  wire sigmoid_table_720_6_sva_dfm_1;
  wire sigmoid_table_721_6_sva_dfm_1;
  wire sigmoid_table_722_6_sva_dfm_1;
  wire sigmoid_table_723_6_sva_dfm_1;
  wire sigmoid_table_724_6_sva_dfm_1;
  wire sigmoid_table_725_6_sva_dfm_1;
  wire sigmoid_table_726_6_sva_dfm_1;
  wire sigmoid_table_727_6_sva_dfm_1;
  wire sigmoid_table_728_6_sva_dfm_1;
  wire sigmoid_table_729_6_sva_dfm_1;
  wire sigmoid_table_730_6_sva_dfm_1;
  wire sigmoid_table_731_6_sva_dfm_1;
  wire sigmoid_table_732_5_sva_dfm_1;
  wire sigmoid_table_733_5_sva_dfm_1;
  wire sigmoid_table_734_5_sva_dfm_1;
  wire sigmoid_table_735_5_sva_dfm_1;
  wire sigmoid_table_736_5_sva_dfm_1;
  wire sigmoid_table_737_5_sva_dfm_1;
  wire sigmoid_table_738_5_sva_dfm_1;
  wire sigmoid_table_739_5_sva_dfm_1;
  wire sigmoid_table_740_5_sva_dfm_1;
  wire sigmoid_table_741_5_sva_dfm_1;
  wire sigmoid_table_742_5_sva_dfm_1;
  wire sigmoid_table_743_5_sva_dfm_1;
  wire sigmoid_table_744_5_sva_dfm_1;
  wire sigmoid_table_745_5_sva_dfm_1;
  wire sigmoid_table_746_5_sva_dfm_1;
  wire sigmoid_table_747_5_sva_dfm_1;
  wire sigmoid_table_748_5_sva_dfm_1;
  wire sigmoid_table_749_5_sva_dfm_1;
  wire sigmoid_table_750_5_sva_dfm_1;
  wire sigmoid_table_751_5_sva_dfm_1;
  wire sigmoid_table_752_5_sva_dfm_1;
  wire sigmoid_table_753_5_sva_dfm_1;
  wire sigmoid_table_754_5_sva_dfm_1;
  wire sigmoid_table_755_5_sva_dfm_1;
  wire sigmoid_table_756_5_sva_dfm_1;
  wire sigmoid_table_757_5_sva_dfm_1;
  wire sigmoid_table_758_5_sva_dfm_1;
  wire sigmoid_table_759_5_sva_dfm_1;
  wire sigmoid_table_760_5_sva_dfm_1;
  wire sigmoid_table_761_5_sva_dfm_1;
  wire sigmoid_table_762_5_sva_dfm_1;
  wire sigmoid_table_763_5_sva_dfm_1;
  wire sigmoid_table_764_5_sva_dfm_1;
  wire sigmoid_table_765_5_sva_dfm_1;
  wire sigmoid_table_766_5_sva_dfm_1;
  wire sigmoid_table_767_5_sva_dfm_1;
  wire sigmoid_table_768_5_sva_dfm_1;
  wire sigmoid_table_769_5_sva_dfm_1;
  wire sigmoid_table_770_5_sva_dfm_1;
  wire sigmoid_table_771_5_sva_dfm_1;
  wire sigmoid_table_772_5_sva_dfm_1;
  wire sigmoid_table_773_5_sva_dfm_1;
  wire sigmoid_table_774_5_sva_dfm_1;
  wire sigmoid_table_775_5_sva_dfm_1;
  wire sigmoid_table_776_5_sva_dfm_1;
  wire sigmoid_table_777_5_sva_dfm_1;
  wire sigmoid_table_778_4_sva_dfm_1;
  wire sigmoid_table_779_4_sva_dfm_1;
  wire sigmoid_table_780_4_sva_dfm_1;
  wire sigmoid_table_781_4_sva_dfm_1;
  wire sigmoid_table_782_4_sva_dfm_1;
  wire sigmoid_table_783_4_sva_dfm_1;
  wire sigmoid_table_784_4_sva_dfm_1;
  wire sigmoid_table_785_4_sva_dfm_1;
  wire sigmoid_table_786_4_sva_dfm_1;
  wire sigmoid_table_787_4_sva_dfm_1;
  wire sigmoid_table_788_4_sva_dfm_1;
  wire sigmoid_table_789_4_sva_dfm_1;
  wire sigmoid_table_790_4_sva_dfm_1;
  wire sigmoid_table_791_4_sva_dfm_1;
  wire sigmoid_table_792_4_sva_dfm_1;
  wire sigmoid_table_793_4_sva_dfm_1;
  wire sigmoid_table_794_4_sva_dfm_1;
  wire sigmoid_table_795_4_sva_dfm_1;
  wire sigmoid_table_796_4_sva_dfm_1;
  wire sigmoid_table_797_4_sva_dfm_1;
  wire sigmoid_table_798_4_sva_dfm_1;
  wire sigmoid_table_799_4_sva_dfm_1;
  wire sigmoid_table_800_4_sva_dfm_1;
  wire sigmoid_table_801_4_sva_dfm_1;
  wire sigmoid_table_802_4_sva_dfm_1;
  wire sigmoid_table_803_4_sva_dfm_1;
  wire sigmoid_table_804_4_sva_dfm_1;
  wire sigmoid_table_805_4_sva_dfm_1;
  wire sigmoid_table_806_4_sva_dfm_1;
  wire sigmoid_table_807_4_sva_dfm_1;
  wire sigmoid_table_808_4_sva_dfm_1;
  wire sigmoid_table_809_4_sva_dfm_1;
  wire sigmoid_table_810_4_sva_dfm_1;
  wire sigmoid_table_811_4_sva_dfm_1;
  wire sigmoid_table_812_4_sva_dfm_1;
  wire sigmoid_table_813_4_sva_dfm_1;
  wire sigmoid_table_814_4_sva_dfm_1;
  wire sigmoid_table_815_4_sva_dfm_1;
  wire sigmoid_table_816_4_sva_dfm_1;
  wire sigmoid_table_817_4_sva_dfm_1;
  wire sigmoid_table_818_4_sva_dfm_1;
  wire sigmoid_table_819_4_sva_dfm_1;
  wire sigmoid_table_820_4_sva_dfm_1;
  wire sigmoid_table_821_4_sva_dfm_1;
  wire sigmoid_table_822_3_sva_dfm_1;
  wire sigmoid_table_823_3_sva_dfm_1;
  wire sigmoid_table_824_3_sva_dfm_1;
  wire sigmoid_table_825_3_sva_dfm_1;
  wire sigmoid_table_826_3_sva_dfm_1;
  wire sigmoid_table_827_3_sva_dfm_1;
  wire sigmoid_table_828_3_sva_dfm_1;
  wire sigmoid_table_829_3_sva_dfm_1;
  wire sigmoid_table_830_3_sva_dfm_1;
  wire sigmoid_table_831_3_sva_dfm_1;
  wire sigmoid_table_832_3_sva_dfm_1;
  wire sigmoid_table_833_3_sva_dfm_1;
  wire sigmoid_table_834_3_sva_dfm_1;
  wire sigmoid_table_835_3_sva_dfm_1;
  wire sigmoid_table_836_3_sva_dfm_1;
  wire sigmoid_table_837_3_sva_dfm_1;
  wire sigmoid_table_838_3_sva_dfm_1;
  wire sigmoid_table_839_3_sva_dfm_1;
  wire sigmoid_table_840_3_sva_dfm_1;
  wire sigmoid_table_841_3_sva_dfm_1;
  wire sigmoid_table_842_3_sva_dfm_1;
  wire sigmoid_table_843_3_sva_dfm_1;
  wire sigmoid_table_844_3_sva_dfm_1;
  wire sigmoid_table_845_3_sva_dfm_1;
  wire sigmoid_table_846_3_sva_dfm_1;
  wire sigmoid_table_847_3_sva_dfm_1;
  wire sigmoid_table_848_3_sva_dfm_1;
  wire sigmoid_table_849_3_sva_dfm_1;
  wire sigmoid_table_850_3_sva_dfm_1;
  wire sigmoid_table_851_3_sva_dfm_1;
  wire sigmoid_table_852_3_sva_dfm_1;
  wire sigmoid_table_853_3_sva_dfm_1;
  wire sigmoid_table_854_3_sva_dfm_1;
  wire sigmoid_table_855_3_sva_dfm_1;
  wire sigmoid_table_856_3_sva_dfm_1;
  wire sigmoid_table_857_3_sva_dfm_1;
  wire sigmoid_table_858_3_sva_dfm_1;
  wire sigmoid_table_859_3_sva_dfm_1;
  wire sigmoid_table_860_3_sva_dfm_1;
  wire sigmoid_table_861_3_sva_dfm_1;
  wire sigmoid_table_862_3_sva_dfm_1;
  wire sigmoid_table_863_3_sva_dfm_1;
  wire sigmoid_table_864_3_sva_dfm_1;
  wire sigmoid_table_865_3_sva_dfm_1;
  wire sigmoid_table_866_3_sva_dfm_1;
  wire sigmoid_table_867_2_sva_dfm_1;
  wire sigmoid_table_868_2_sva_dfm_1;
  wire sigmoid_table_869_2_sva_dfm_1;
  wire sigmoid_table_870_2_sva_dfm_1;
  wire sigmoid_table_871_2_sva_dfm_1;
  wire sigmoid_table_872_2_sva_dfm_1;
  wire sigmoid_table_873_2_sva_dfm_1;
  wire sigmoid_table_874_2_sva_dfm_1;
  wire sigmoid_table_875_2_sva_dfm_1;
  wire sigmoid_table_876_2_sva_dfm_1;
  wire sigmoid_table_877_2_sva_dfm_1;
  wire sigmoid_table_878_2_sva_dfm_1;
  wire sigmoid_table_879_2_sva_dfm_1;
  wire sigmoid_table_880_2_sva_dfm_1;
  wire sigmoid_table_881_2_sva_dfm_1;
  wire sigmoid_table_882_2_sva_dfm_1;
  wire sigmoid_table_883_2_sva_dfm_1;
  wire sigmoid_table_884_2_sva_dfm_1;
  wire sigmoid_table_885_2_sva_dfm_1;
  wire sigmoid_table_886_2_sva_dfm_1;
  wire sigmoid_table_887_2_sva_dfm_1;
  wire sigmoid_table_888_2_sva_dfm_1;
  wire sigmoid_table_889_2_sva_dfm_1;
  wire sigmoid_table_890_2_sva_dfm_1;
  wire sigmoid_table_891_2_sva_dfm_1;
  wire sigmoid_table_892_2_sva_dfm_1;
  wire sigmoid_table_893_2_sva_dfm_1;
  wire sigmoid_table_894_2_sva_dfm_1;
  wire sigmoid_table_895_2_sva_dfm_1;
  wire sigmoid_table_896_2_sva_dfm_1;
  wire sigmoid_table_897_2_sva_dfm_1;
  wire sigmoid_table_898_2_sva_dfm_1;
  wire sigmoid_table_899_2_sva_dfm_1;
  wire sigmoid_table_900_2_sva_dfm_1;
  wire sigmoid_table_901_2_sva_dfm_1;
  wire sigmoid_table_902_2_sva_dfm_1;
  wire sigmoid_table_903_2_sva_dfm_1;
  wire sigmoid_table_904_2_sva_dfm_1;
  wire sigmoid_table_905_2_sva_dfm_1;
  wire sigmoid_table_906_2_sva_dfm_1;
  wire sigmoid_table_907_2_sva_dfm_1;
  wire sigmoid_table_908_2_sva_dfm_1;
  wire sigmoid_table_909_2_sva_dfm_1;
  wire sigmoid_table_910_2_sva_dfm_1;
  wire sigmoid_table_911_1_sva_dfm_1;
  wire sigmoid_table_912_1_sva_dfm_1;
  wire sigmoid_table_913_1_sva_dfm_1;
  wire sigmoid_table_914_1_sva_dfm_1;
  wire sigmoid_table_915_1_sva_dfm_1;
  wire sigmoid_table_916_1_sva_dfm_1;
  wire sigmoid_table_917_1_sva_dfm_1;
  wire sigmoid_table_918_1_sva_dfm_1;
  wire sigmoid_table_919_1_sva_dfm_1;
  wire sigmoid_table_920_1_sva_dfm_1;
  wire sigmoid_table_921_1_sva_dfm_1;
  wire sigmoid_table_922_1_sva_dfm_1;
  wire sigmoid_table_923_1_sva_dfm_1;
  wire sigmoid_table_924_1_sva_dfm_1;
  wire sigmoid_table_925_1_sva_dfm_1;
  wire sigmoid_table_926_1_sva_dfm_1;
  wire sigmoid_table_927_1_sva_dfm_1;
  wire sigmoid_table_928_1_sva_dfm_1;
  wire sigmoid_table_929_1_sva_dfm_1;
  wire sigmoid_table_930_1_sva_dfm_1;
  wire sigmoid_table_931_1_sva_dfm_1;
  wire sigmoid_table_932_1_sva_dfm_1;
  wire sigmoid_table_933_1_sva_dfm_1;
  wire sigmoid_table_934_1_sva_dfm_1;
  wire sigmoid_table_935_1_sva_dfm_1;
  wire sigmoid_table_936_1_sva_dfm_1;
  wire sigmoid_table_937_1_sva_dfm_1;
  wire sigmoid_table_938_1_sva_dfm_1;
  wire sigmoid_table_939_1_sva_dfm_1;
  wire sigmoid_table_940_1_sva_dfm_1;
  wire sigmoid_table_941_1_sva_dfm_1;
  wire sigmoid_table_942_1_sva_dfm_1;
  wire sigmoid_table_943_1_sva_dfm_1;
  wire sigmoid_table_944_1_sva_dfm_1;
  wire sigmoid_table_945_1_sva_dfm_1;
  wire sigmoid_table_946_1_sva_dfm_1;
  wire sigmoid_table_947_1_sva_dfm_1;
  wire sigmoid_table_948_1_sva_dfm_1;
  wire sigmoid_table_949_1_sva_dfm_1;
  wire sigmoid_table_950_1_sva_dfm_1;
  wire sigmoid_table_951_1_sva_dfm_1;
  wire sigmoid_table_952_1_sva_dfm_1;
  wire sigmoid_table_953_1_sva_dfm_1;
  wire sigmoid_table_954_1_sva_dfm_1;
  wire sigmoid_table_113_1_sva_dfm_1;
  wire sigmoid_table_114_1_sva_dfm_1;
  wire sigmoid_table_115_1_sva_dfm_1;
  wire sigmoid_table_116_1_sva_dfm_1;
  wire sigmoid_table_117_1_sva_dfm_1;
  wire sigmoid_table_118_1_sva_dfm_1;
  wire sigmoid_table_119_1_sva_dfm_1;
  wire sigmoid_table_120_1_sva_dfm_1;
  wire sigmoid_table_121_1_sva_dfm_1;
  wire sigmoid_table_122_1_sva_dfm_1;
  wire sigmoid_table_123_1_sva_dfm_1;
  wire sigmoid_table_124_1_sva_dfm_1;
  wire sigmoid_table_125_1_sva_dfm_1;
  wire sigmoid_table_126_1_sva_dfm_1;
  wire sigmoid_table_127_1_sva_dfm_1;
  wire sigmoid_table_128_1_sva_dfm_1;
  wire sigmoid_table_129_1_sva_dfm_1;
  wire sigmoid_table_130_1_sva_dfm_1;
  wire sigmoid_table_131_1_sva_dfm_1;
  wire sigmoid_table_132_1_sva_dfm_1;
  wire sigmoid_table_133_1_sva_dfm_1;
  wire sigmoid_table_134_1_sva_dfm_1;
  wire sigmoid_table_135_1_sva_dfm_1;
  wire sigmoid_table_136_1_sva_dfm_1;
  wire sigmoid_table_137_1_sva_dfm_1;
  wire sigmoid_table_138_1_sva_dfm_1;
  wire sigmoid_table_184_1_sva_dfm_1;
  wire sigmoid_table_185_1_sva_dfm_1;
  wire sigmoid_table_186_1_sva_dfm_1;
  wire sigmoid_table_187_1_sva_dfm_1;
  wire sigmoid_table_188_1_sva_dfm_1;
  wire sigmoid_table_189_1_sva_dfm_1;
  wire sigmoid_table_190_1_sva_dfm_1;
  wire sigmoid_table_191_1_sva_dfm_1;
  wire sigmoid_table_192_1_sva_dfm_1;
  wire sigmoid_table_193_1_sva_dfm_1;
  wire sigmoid_table_217_1_sva_dfm_1;
  wire sigmoid_table_218_1_sva_dfm_1;
  wire sigmoid_table_219_1_sva_dfm_1;
  wire sigmoid_table_220_1_sva_dfm_1;
  wire sigmoid_table_221_1_sva_dfm_1;
  wire sigmoid_table_222_1_sva_dfm_1;
  wire sigmoid_table_239_1_sva_dfm_1;
  wire sigmoid_table_240_1_sva_dfm_1;
  wire sigmoid_table_241_1_sva_dfm_1;
  wire sigmoid_table_242_1_sva_dfm_1;
  wire sigmoid_table_255_1_sva_dfm_1;
  wire sigmoid_table_256_1_sva_dfm_1;
  wire sigmoid_table_257_1_sva_dfm_1;
  wire sigmoid_table_258_1_sva_dfm_1;
  wire sigmoid_table_268_1_sva_dfm_1;
  wire sigmoid_table_269_1_sva_dfm_1;
  wire sigmoid_table_270_1_sva_dfm_1;
  wire sigmoid_table_279_1_sva_dfm_1;
  wire sigmoid_table_280_1_sva_dfm_1;
  wire sigmoid_table_281_1_sva_dfm_1;
  wire sigmoid_table_288_1_sva_dfm_1;
  wire sigmoid_table_289_1_sva_dfm_1;
  wire sigmoid_table_290_1_sva_dfm_1;
  wire sigmoid_table_297_1_sva_dfm_1;
  wire sigmoid_table_298_1_sva_dfm_1;
  wire sigmoid_table_304_1_sva_dfm_1;
  wire sigmoid_table_305_1_sva_dfm_1;
  wire sigmoid_table_311_1_sva_dfm_1;
  wire sigmoid_table_317_1_sva_dfm_1;
  wire sigmoid_table_322_1_sva_dfm_1;
  wire sigmoid_table_323_1_sva_dfm_1;
  wire sigmoid_table_328_1_sva_dfm_1;
  wire sigmoid_table_332_1_sva_dfm_1;
  wire sigmoid_table_333_1_sva_dfm_1;
  wire sigmoid_table_337_1_sva_dfm_1;
  wire sigmoid_table_341_1_sva_dfm_1;
  wire sigmoid_table_345_1_sva_dfm_1;
  wire sigmoid_table_349_1_sva_dfm_1;
  wire sigmoid_table_353_1_sva_dfm_1;
  wire sigmoid_table_356_1_sva_dfm_1;
  wire sigmoid_table_363_1_sva_dfm_1;
  wire sigmoid_table_366_1_sva_dfm_1;
  wire sigmoid_table_374_1_sva_dfm_1;
  wire sigmoid_table_377_1_sva_dfm_1;
  wire sigmoid_table_382_1_sva_dfm_1;
  wire sigmoid_table_384_1_sva_dfm_1;
  wire sigmoid_table_389_1_sva_dfm_1;
  wire sigmoid_table_391_1_sva_dfm_1;
  wire sigmoid_table_393_1_sva_dfm_1;
  wire sigmoid_table_407_1_sva_dfm_1;
  wire sigmoid_table_409_1_sva_dfm_1;
  wire sigmoid_table_414_1_sva_dfm_1;
  wire sigmoid_table_416_1_sva_dfm_1;
  wire sigmoid_table_419_1_sva_dfm_1;
  wire sigmoid_table_424_1_sva_dfm_1;
  wire sigmoid_table_427_1_sva_dfm_1;
  wire sigmoid_table_430_1_sva_dfm_1;
  wire sigmoid_table_433_1_sva_dfm_1;
  wire sigmoid_table_437_1_sva_dfm_1;
  wire sigmoid_table_440_1_sva_dfm_1;
  wire sigmoid_table_444_1_sva_dfm_1;
  wire sigmoid_table_445_1_sva_dfm_1;
  wire sigmoid_table_449_1_sva_dfm_1;
  wire sigmoid_table_454_1_sva_dfm_1;
  wire sigmoid_table_460_1_sva_dfm_1;
  wire sigmoid_table_461_1_sva_dfm_1;
  wire sigmoid_table_468_1_sva_dfm_1;
  wire sigmoid_table_469_1_sva_dfm_1;
  wire sigmoid_table_479_1_sva_dfm_1;
  wire sigmoid_table_480_1_sva_dfm_1;
  wire sigmoid_table_481_1_sva_dfm_1;
  wire sigmoid_table_482_1_sva_dfm_1;
  wire sigmoid_table_536_1_sva_dfm_1;
  wire sigmoid_table_537_1_sva_dfm_1;
  wire sigmoid_table_538_1_sva_dfm_1;
  wire sigmoid_table_539_1_sva_dfm_1;
  wire sigmoid_table_540_1_sva_dfm_1;
  wire sigmoid_table_541_1_sva_dfm_1;
  wire sigmoid_table_552_1_sva_dfm_1;
  wire sigmoid_table_553_1_sva_dfm_1;
  wire sigmoid_table_554_1_sva_dfm_1;
  wire sigmoid_table_561_1_sva_dfm_1;
  wire sigmoid_table_562_1_sva_dfm_1;
  wire sigmoid_table_568_1_sva_dfm_1;
  wire sigmoid_table_569_1_sva_dfm_1;
  wire sigmoid_table_574_1_sva_dfm_1;
  wire sigmoid_table_578_1_sva_dfm_1;
  wire sigmoid_table_583_1_sva_dfm_1;
  wire sigmoid_table_586_1_sva_dfm_1;
  wire sigmoid_table_590_1_sva_dfm_1;
  wire sigmoid_table_593_1_sva_dfm_1;
  wire sigmoid_table_596_1_sva_dfm_1;
  wire sigmoid_table_599_1_sva_dfm_1;
  wire sigmoid_table_602_1_sva_dfm_1;
  wire sigmoid_table_607_1_sva_dfm_1;
  wire sigmoid_table_612_1_sva_dfm_1;
  wire sigmoid_table_619_1_sva_dfm_1;
  wire sigmoid_table_621_1_sva_dfm_1;
  wire sigmoid_table_623_1_sva_dfm_1;
  wire sigmoid_table_625_1_sva_dfm_1;
  wire sigmoid_table_627_1_sva_dfm_1;
  wire sigmoid_table_629_1_sva_dfm_1;
  wire sigmoid_table_638_1_sva_dfm_1;
  wire sigmoid_table_643_1_sva_dfm_1;
  wire sigmoid_table_645_1_sva_dfm_1;
  wire sigmoid_table_648_1_sva_dfm_1;
  wire sigmoid_table_653_1_sva_dfm_1;
  wire sigmoid_table_656_1_sva_dfm_1;
  wire sigmoid_table_659_1_sva_dfm_1;
  wire sigmoid_table_662_1_sva_dfm_1;
  wire sigmoid_table_665_1_sva_dfm_1;
  wire sigmoid_table_669_1_sva_dfm_1;
  wire sigmoid_table_672_1_sva_dfm_1;
  wire sigmoid_table_676_1_sva_dfm_1;
  wire sigmoid_table_680_1_sva_dfm_1;
  wire sigmoid_table_684_1_sva_dfm_1;
  wire sigmoid_table_688_1_sva_dfm_1;
  wire sigmoid_table_693_1_sva_dfm_1;
  wire sigmoid_table_697_1_sva_dfm_1;
  wire sigmoid_table_698_1_sva_dfm_1;
  wire sigmoid_table_703_1_sva_dfm_1;
  wire sigmoid_table_708_1_sva_dfm_1;
  wire sigmoid_table_709_1_sva_dfm_1;
  wire sigmoid_table_714_1_sva_dfm_1;
  wire sigmoid_table_715_1_sva_dfm_1;
  wire sigmoid_table_721_1_sva_dfm_1;
  wire sigmoid_table_722_1_sva_dfm_1;
  wire sigmoid_table_728_1_sva_dfm_1;
  wire sigmoid_table_729_1_sva_dfm_1;
  wire sigmoid_table_737_1_sva_dfm_1;
  wire sigmoid_table_738_1_sva_dfm_1;
  wire sigmoid_table_746_1_sva_dfm_1;
  wire sigmoid_table_747_1_sva_dfm_1;
  wire sigmoid_table_757_1_sva_dfm_1;
  wire sigmoid_table_758_1_sva_dfm_1;
  wire sigmoid_table_759_1_sva_dfm_1;
  wire sigmoid_table_770_1_sva_dfm_1;
  wire sigmoid_table_771_1_sva_dfm_1;
  wire sigmoid_table_772_1_sva_dfm_1;
  wire sigmoid_table_773_1_sva_dfm_1;
  wire sigmoid_table_786_1_sva_dfm_1;
  wire sigmoid_table_787_1_sva_dfm_1;
  wire sigmoid_table_788_1_sva_dfm_1;
  wire sigmoid_table_789_1_sva_dfm_1;
  wire sigmoid_table_790_1_sva_dfm_1;
  wire sigmoid_table_808_1_sva_dfm_1;
  wire sigmoid_table_809_1_sva_dfm_1;
  wire sigmoid_table_810_1_sva_dfm_1;
  wire sigmoid_table_811_1_sva_dfm_1;
  wire sigmoid_table_812_1_sva_dfm_1;
  wire sigmoid_table_813_1_sva_dfm_1;
  wire sigmoid_table_814_1_sva_dfm_1;
  wire sigmoid_table_841_1_sva_dfm_1;
  wire sigmoid_table_842_1_sva_dfm_1;
  wire sigmoid_table_843_1_sva_dfm_1;
  wire sigmoid_table_844_1_sva_dfm_1;
  wire sigmoid_table_845_1_sva_dfm_1;
  wire sigmoid_table_846_1_sva_dfm_1;
  wire sigmoid_table_847_1_sva_dfm_1;
  wire sigmoid_table_848_1_sva_dfm_1;
  wire sigmoid_table_849_1_sva_dfm_1;
  wire sigmoid_table_850_1_sva_dfm_1;
  wire sigmoid_table_851_1_sva_dfm_1;
  wire sigmoid_table_852_1_sva_dfm_1;
  wire sigmoid_table_442_8_sva_dfm_1;
  wire sigmoid_table_443_8_sva_dfm_1;
  wire sigmoid_table_444_8_sva_dfm_1;
  wire sigmoid_table_445_8_sva_dfm_1;
  wire sigmoid_table_446_8_sva_dfm_1;
  wire sigmoid_table_447_8_sva_dfm_1;
  wire sigmoid_table_448_8_sva_dfm_1;
  wire sigmoid_table_449_8_sva_dfm_1;
  wire sigmoid_table_450_8_sva_dfm_1;
  wire sigmoid_table_451_8_sva_dfm_1;
  wire sigmoid_table_452_8_sva_dfm_1;
  wire sigmoid_table_453_8_sva_dfm_1;
  wire sigmoid_table_454_8_sva_dfm_1;
  wire sigmoid_table_455_8_sva_dfm_1;
  wire sigmoid_table_456_8_sva_dfm_1;
  wire sigmoid_table_457_8_sva_dfm_1;
  wire sigmoid_table_458_8_sva_dfm_1;
  wire sigmoid_table_459_8_sva_dfm_1;
  wire sigmoid_table_460_8_sva_dfm_1;
  wire sigmoid_table_461_8_sva_dfm_1;
  wire sigmoid_table_462_8_sva_dfm_1;
  wire sigmoid_table_463_8_sva_dfm_1;
  wire sigmoid_table_464_8_sva_dfm_1;
  wire sigmoid_table_465_8_sva_dfm_1;
  wire sigmoid_table_466_8_sva_dfm_1;
  wire sigmoid_table_467_8_sva_dfm_1;
  wire sigmoid_table_468_8_sva_dfm_1;
  wire sigmoid_table_469_8_sva_dfm_1;
  wire sigmoid_table_470_8_sva_dfm_1;
  wire sigmoid_table_471_8_sva_dfm_1;
  wire sigmoid_table_472_8_sva_dfm_1;
  wire sigmoid_table_473_8_sva_dfm_1;
  wire sigmoid_table_474_8_sva_dfm_1;
  wire sigmoid_table_475_8_sva_dfm_1;
  wire sigmoid_table_476_8_sva_dfm_1;
  wire sigmoid_table_477_8_sva_dfm_1;
  wire sigmoid_table_478_8_sva_dfm_1;
  wire sigmoid_table_479_8_sva_dfm_1;
  wire sigmoid_table_480_7_sva_dfm_1;
  wire sigmoid_table_481_7_sva_dfm_1;
  wire sigmoid_table_482_7_sva_dfm_1;
  wire sigmoid_table_483_7_sva_dfm_1;
  wire sigmoid_table_484_7_sva_dfm_1;
  wire sigmoid_table_485_7_sva_dfm_1;
  wire sigmoid_table_486_7_sva_dfm_1;
  wire sigmoid_table_487_7_sva_dfm_1;
  wire sigmoid_table_488_7_sva_dfm_1;
  wire sigmoid_table_489_7_sva_dfm_1;
  wire sigmoid_table_490_7_sva_dfm_1;
  wire sigmoid_table_491_7_sva_dfm_1;
  wire sigmoid_table_492_7_sva_dfm_1;
  wire sigmoid_table_493_7_sva_dfm_1;
  wire sigmoid_table_494_7_sva_dfm_1;
  wire sigmoid_table_495_7_sva_dfm_1;
  wire sigmoid_table_496_6_sva_dfm_1;
  wire sigmoid_table_497_6_sva_dfm_1;
  wire sigmoid_table_498_6_sva_dfm_1;
  wire sigmoid_table_499_6_sva_dfm_1;
  wire sigmoid_table_500_6_sva_dfm_1;
  wire sigmoid_table_501_6_sva_dfm_1;
  wire sigmoid_table_502_6_sva_dfm_1;
  wire sigmoid_table_503_6_sva_dfm_1;
  wire sigmoid_table_504_5_sva_dfm_1;
  wire sigmoid_table_505_5_sva_dfm_1;
  wire sigmoid_table_506_5_sva_dfm_1;
  wire sigmoid_table_507_5_sva_dfm_1;
  wire sigmoid_table_508_4_sva_dfm_1;
  wire sigmoid_table_509_4_sva_dfm_1;
  wire sigmoid_table_510_3_sva_dfm_1;
  wire sigmoid_table_511_2_sva_dfm_1;
  wire sigmoid_table_158_2_sva_dfm_1;
  wire sigmoid_table_159_2_sva_dfm_1;
  wire sigmoid_table_160_2_sva_dfm_1;
  wire sigmoid_table_161_2_sva_dfm_1;
  wire sigmoid_table_162_2_sva_dfm_1;
  wire sigmoid_table_163_2_sva_dfm_1;
  wire sigmoid_table_164_2_sva_dfm_1;
  wire sigmoid_table_165_2_sva_dfm_1;
  wire sigmoid_table_166_2_sva_dfm_1;
  wire sigmoid_table_167_2_sva_dfm_1;
  wire sigmoid_table_168_2_sva_dfm_1;
  wire sigmoid_table_169_2_sva_dfm_1;
  wire sigmoid_table_170_2_sva_dfm_1;
  wire sigmoid_table_171_2_sva_dfm_1;
  wire sigmoid_table_172_2_sva_dfm_1;
  wire sigmoid_table_173_2_sva_dfm_1;
  wire sigmoid_table_174_2_sva_dfm_1;
  wire sigmoid_table_175_2_sva_dfm_1;
  wire sigmoid_table_176_2_sva_dfm_1;
  wire sigmoid_table_177_2_sva_dfm_1;
  wire sigmoid_table_178_2_sva_dfm_1;
  wire sigmoid_table_179_2_sva_dfm_1;
  wire sigmoid_table_180_2_sva_dfm_1;
  wire sigmoid_table_181_2_sva_dfm_1;
  wire sigmoid_table_182_2_sva_dfm_1;
  wire sigmoid_table_183_2_sva_dfm_1;
  wire sigmoid_table_229_2_sva_dfm_1;
  wire sigmoid_table_230_2_sva_dfm_1;
  wire sigmoid_table_231_2_sva_dfm_1;
  wire sigmoid_table_232_2_sva_dfm_1;
  wire sigmoid_table_233_2_sva_dfm_1;
  wire sigmoid_table_234_2_sva_dfm_1;
  wire sigmoid_table_235_2_sva_dfm_1;
  wire sigmoid_table_236_2_sva_dfm_1;
  wire sigmoid_table_237_2_sva_dfm_1;
  wire sigmoid_table_238_2_sva_dfm_1;
  wire sigmoid_table_262_2_sva_dfm_1;
  wire sigmoid_table_263_2_sva_dfm_1;
  wire sigmoid_table_264_2_sva_dfm_1;
  wire sigmoid_table_265_2_sva_dfm_1;
  wire sigmoid_table_266_2_sva_dfm_1;
  wire sigmoid_table_267_2_sva_dfm_1;
  wire sigmoid_table_284_2_sva_dfm_1;
  wire sigmoid_table_285_2_sva_dfm_1;
  wire sigmoid_table_286_2_sva_dfm_1;
  wire sigmoid_table_287_2_sva_dfm_1;
  wire sigmoid_table_301_2_sva_dfm_1;
  wire sigmoid_table_302_2_sva_dfm_1;
  wire sigmoid_table_303_2_sva_dfm_1;
  wire sigmoid_table_314_2_sva_dfm_1;
  wire sigmoid_table_315_2_sva_dfm_1;
  wire sigmoid_table_316_2_sva_dfm_1;
  wire sigmoid_table_325_2_sva_dfm_1;
  wire sigmoid_table_326_2_sva_dfm_1;
  wire sigmoid_table_327_2_sva_dfm_1;
  wire sigmoid_table_335_2_sva_dfm_1;
  wire sigmoid_table_336_2_sva_dfm_1;
  wire sigmoid_table_343_2_sva_dfm_1;
  wire sigmoid_table_344_2_sva_dfm_1;
  wire sigmoid_table_351_2_sva_dfm_1;
  wire sigmoid_table_352_2_sva_dfm_1;
  wire sigmoid_table_358_2_sva_dfm_1;
  wire sigmoid_table_359_2_sva_dfm_1;
  wire sigmoid_table_364_2_sva_dfm_1;
  wire sigmoid_table_365_2_sva_dfm_1;
  wire sigmoid_table_370_2_sva_dfm_1;
  wire sigmoid_table_371_2_sva_dfm_1;
  wire sigmoid_table_376_2_sva_dfm_1;
  wire sigmoid_table_381_2_sva_dfm_1;
  wire sigmoid_table_386_2_sva_dfm_1;
  wire sigmoid_table_390_2_sva_dfm_1;
  wire sigmoid_table_395_2_sva_dfm_1;
  wire sigmoid_table_399_2_sva_dfm_1;
  wire sigmoid_table_403_2_sva_dfm_1;
  wire sigmoid_table_406_2_sva_dfm_1;
  wire sigmoid_table_410_2_sva_dfm_1;
  wire sigmoid_table_417_2_sva_dfm_1;
  wire sigmoid_table_420_2_sva_dfm_1;
  wire sigmoid_table_423_2_sva_dfm_1;
  wire sigmoid_table_432_2_sva_dfm_1;
  wire sigmoid_table_435_2_sva_dfm_1;
  wire sigmoid_table_438_2_sva_dfm_1;
  wire sigmoid_table_441_2_sva_dfm_1;
  wire sigmoid_table_446_2_sva_dfm_1;
  wire sigmoid_table_451_2_sva_dfm_1;
  wire sigmoid_table_456_2_sva_dfm_1;
  wire sigmoid_table_463_2_sva_dfm_1;
  wire sigmoid_table_465_2_sva_dfm_1;
  wire sigmoid_table_470_2_sva_dfm_1;
  wire sigmoid_table_472_2_sva_dfm_1;
  wire sigmoid_table_474_2_sva_dfm_1;
  wire sigmoid_table_483_2_sva_dfm_1;
  wire sigmoid_table_485_2_sva_dfm_1;
  wire sigmoid_table_487_2_sva_dfm_1;
  wire sigmoid_table_489_2_sva_dfm_1;
  wire sigmoid_table_491_2_sva_dfm_1;
  wire sigmoid_table_493_2_sva_dfm_1;
  wire sigmoid_table_495_2_sva_dfm_1;
  wire sigmoid_table_497_2_sva_dfm_1;
  wire sigmoid_table_499_2_sva_dfm_1;
  wire sigmoid_table_501_2_sva_dfm_1;
  wire sigmoid_table_503_2_sva_dfm_1;
  wire sigmoid_table_505_2_sva_dfm_1;
  wire sigmoid_table_507_2_sva_dfm_1;
  wire sigmoid_table_509_2_sva_dfm_1;
  wire sigmoid_table_513_2_sva_dfm_1;
  wire sigmoid_table_515_2_sva_dfm_1;
  wire sigmoid_table_542_2_sva_dfm_1;
  wire sigmoid_table_544_2_sva_dfm_1;
  wire sigmoid_table_546_2_sva_dfm_1;
  wire sigmoid_table_548_2_sva_dfm_1;
  wire sigmoid_table_555_2_sva_dfm_1;
  wire sigmoid_table_557_2_sva_dfm_1;
  wire sigmoid_table_564_2_sva_dfm_1;
  wire sigmoid_table_566_2_sva_dfm_1;
  wire sigmoid_table_571_2_sva_dfm_1;
  wire sigmoid_table_576_2_sva_dfm_1;
  wire sigmoid_table_579_2_sva_dfm_1;
  wire sigmoid_table_581_2_sva_dfm_1;
  wire sigmoid_table_584_2_sva_dfm_1;
  wire sigmoid_table_587_2_sva_dfm_1;
  wire sigmoid_table_595_2_sva_dfm_1;
  wire sigmoid_table_598_2_sva_dfm_1;
  wire sigmoid_table_605_2_sva_dfm_1;
  wire sigmoid_table_608_2_sva_dfm_1;
  wire sigmoid_table_611_2_sva_dfm_1;
  wire sigmoid_table_615_2_sva_dfm_1;
  wire sigmoid_table_622_2_sva_dfm_1;
  wire sigmoid_table_626_2_sva_dfm_1;
  wire sigmoid_table_630_2_sva_dfm_1;
  wire sigmoid_table_631_2_sva_dfm_1;
  wire sigmoid_table_635_2_sva_dfm_1;
  wire sigmoid_table_639_2_sva_dfm_1;
  wire sigmoid_table_640_2_sva_dfm_1;
  wire sigmoid_table_644_2_sva_dfm_1;
  wire sigmoid_table_649_2_sva_dfm_1;
  wire sigmoid_table_650_2_sva_dfm_1;
  wire sigmoid_table_655_2_sva_dfm_1;
  wire sigmoid_table_661_2_sva_dfm_1;
  wire sigmoid_table_667_2_sva_dfm_1;
  wire sigmoid_table_668_2_sva_dfm_1;
  wire sigmoid_table_674_2_sva_dfm_1;
  wire sigmoid_table_675_2_sva_dfm_1;
  wire sigmoid_table_682_2_sva_dfm_1;
  wire sigmoid_table_683_2_sva_dfm_1;
  wire sigmoid_table_690_2_sva_dfm_1;
  wire sigmoid_table_691_2_sva_dfm_1;
  wire sigmoid_table_692_2_sva_dfm_1;
  wire sigmoid_table_700_2_sva_dfm_1;
  wire sigmoid_table_701_2_sva_dfm_1;
  wire sigmoid_table_702_2_sva_dfm_1;
  wire sigmoid_table_711_2_sva_dfm_1;
  wire sigmoid_table_712_2_sva_dfm_1;
  wire sigmoid_table_713_2_sva_dfm_1;
  wire sigmoid_table_724_2_sva_dfm_1;
  wire sigmoid_table_725_2_sva_dfm_1;
  wire sigmoid_table_726_2_sva_dfm_1;
  wire sigmoid_table_727_2_sva_dfm_1;
  wire sigmoid_table_741_2_sva_dfm_1;
  wire sigmoid_table_742_2_sva_dfm_1;
  wire sigmoid_table_743_2_sva_dfm_1;
  wire sigmoid_table_744_2_sva_dfm_1;
  wire sigmoid_table_745_2_sva_dfm_1;
  wire sigmoid_table_763_2_sva_dfm_1;
  wire sigmoid_table_764_2_sva_dfm_1;
  wire sigmoid_table_765_2_sva_dfm_1;
  wire sigmoid_table_766_2_sva_dfm_1;
  wire sigmoid_table_767_2_sva_dfm_1;
  wire sigmoid_table_768_2_sva_dfm_1;
  wire sigmoid_table_769_2_sva_dfm_1;
  wire sigmoid_table_796_2_sva_dfm_1;
  wire sigmoid_table_797_2_sva_dfm_1;
  wire sigmoid_table_798_2_sva_dfm_1;
  wire sigmoid_table_799_2_sva_dfm_1;
  wire sigmoid_table_800_2_sva_dfm_1;
  wire sigmoid_table_801_2_sva_dfm_1;
  wire sigmoid_table_802_2_sva_dfm_1;
  wire sigmoid_table_803_2_sva_dfm_1;
  wire sigmoid_table_804_2_sva_dfm_1;
  wire sigmoid_table_805_2_sva_dfm_1;
  wire sigmoid_table_806_2_sva_dfm_1;
  wire sigmoid_table_807_2_sva_dfm_1;
  wire sigmoid_table_388_7_sva_dfm_1;
  wire sigmoid_table_389_7_sva_dfm_1;
  wire sigmoid_table_390_7_sva_dfm_1;
  wire sigmoid_table_391_7_sva_dfm_1;
  wire sigmoid_table_392_7_sva_dfm_1;
  wire sigmoid_table_393_7_sva_dfm_1;
  wire sigmoid_table_394_7_sva_dfm_1;
  wire sigmoid_table_395_7_sva_dfm_1;
  wire sigmoid_table_396_7_sva_dfm_1;
  wire sigmoid_table_397_7_sva_dfm_1;
  wire sigmoid_table_398_7_sva_dfm_1;
  wire sigmoid_table_399_7_sva_dfm_1;
  wire sigmoid_table_400_7_sva_dfm_1;
  wire sigmoid_table_401_7_sva_dfm_1;
  wire sigmoid_table_402_7_sva_dfm_1;
  wire sigmoid_table_403_7_sva_dfm_1;
  wire sigmoid_table_404_7_sva_dfm_1;
  wire sigmoid_table_405_7_sva_dfm_1;
  wire sigmoid_table_406_7_sva_dfm_1;
  wire sigmoid_table_407_7_sva_dfm_1;
  wire sigmoid_table_408_7_sva_dfm_1;
  wire sigmoid_table_409_7_sva_dfm_1;
  wire sigmoid_table_410_7_sva_dfm_1;
  wire sigmoid_table_411_7_sva_dfm_1;
  wire sigmoid_table_412_7_sva_dfm_1;
  wire sigmoid_table_413_7_sva_dfm_1;
  wire sigmoid_table_414_7_sva_dfm_1;
  wire sigmoid_table_415_7_sva_dfm_1;
  wire sigmoid_table_416_7_sva_dfm_1;
  wire sigmoid_table_417_7_sva_dfm_1;
  wire sigmoid_table_418_7_sva_dfm_1;
  wire sigmoid_table_419_6_sva_dfm_1;
  wire sigmoid_table_420_6_sva_dfm_1;
  wire sigmoid_table_421_6_sva_dfm_1;
  wire sigmoid_table_422_6_sva_dfm_1;
  wire sigmoid_table_423_6_sva_dfm_1;
  wire sigmoid_table_424_6_sva_dfm_1;
  wire sigmoid_table_425_6_sva_dfm_1;
  wire sigmoid_table_426_6_sva_dfm_1;
  wire sigmoid_table_427_6_sva_dfm_1;
  wire sigmoid_table_428_6_sva_dfm_1;
  wire sigmoid_table_429_6_sva_dfm_1;
  wire sigmoid_table_430_6_sva_dfm_1;
  wire sigmoid_table_431_5_sva_dfm_1;
  wire sigmoid_table_432_5_sva_dfm_1;
  wire sigmoid_table_433_5_sva_dfm_1;
  wire sigmoid_table_434_5_sva_dfm_1;
  wire sigmoid_table_435_5_sva_dfm_1;
  wire sigmoid_table_436_5_sva_dfm_1;
  wire sigmoid_table_437_4_sva_dfm_1;
  wire sigmoid_table_438_4_sva_dfm_1;
  wire sigmoid_table_439_3_sva_dfm_1;
  wire sigmoid_table_440_3_sva_dfm_1;
  wire sigmoid_table_545_7_sva_dfm_1;
  wire sigmoid_table_546_7_sva_dfm_1;
  wire sigmoid_table_547_7_sva_dfm_1;
  wire sigmoid_table_548_7_sva_dfm_1;
  wire sigmoid_table_549_7_sva_dfm_1;
  wire sigmoid_table_550_7_sva_dfm_1;
  wire sigmoid_table_551_7_sva_dfm_1;
  wire sigmoid_table_552_7_sva_dfm_1;
  wire sigmoid_table_553_7_sva_dfm_1;
  wire sigmoid_table_554_7_sva_dfm_1;
  wire sigmoid_table_555_7_sva_dfm_1;
  wire sigmoid_table_556_7_sva_dfm_1;
  wire sigmoid_table_557_7_sva_dfm_1;
  wire sigmoid_table_558_7_sva_dfm_1;
  wire sigmoid_table_559_7_sva_dfm_1;
  wire sigmoid_table_560_7_sva_dfm_1;
  wire sigmoid_table_561_7_sva_dfm_1;
  wire sigmoid_table_562_7_sva_dfm_1;
  wire sigmoid_table_563_6_sva_dfm_1;
  wire sigmoid_table_564_6_sva_dfm_1;
  wire sigmoid_table_565_6_sva_dfm_1;
  wire sigmoid_table_566_6_sva_dfm_1;
  wire sigmoid_table_567_6_sva_dfm_1;
  wire sigmoid_table_568_6_sva_dfm_1;
  wire sigmoid_table_569_6_sva_dfm_1;
  wire sigmoid_table_570_6_sva_dfm_1;
  wire sigmoid_table_571_6_sva_dfm_1;
  wire sigmoid_table_572_6_sva_dfm_1;
  wire sigmoid_table_573_5_sva_dfm_1;
  wire sigmoid_table_574_5_sva_dfm_1;
  wire sigmoid_table_575_5_sva_dfm_1;
  wire sigmoid_table_576_5_sva_dfm_1;
  wire sigmoid_table_577_5_sva_dfm_1;
  wire sigmoid_table_578_4_sva_dfm_1;
  wire sigmoid_table_579_4_sva_dfm_1;
  wire sigmoid_table_580_3_sva_dfm_1;
  wire sigmoid_table_202_3_sva_dfm_1;
  wire sigmoid_table_203_3_sva_dfm_1;
  wire sigmoid_table_204_3_sva_dfm_1;
  wire sigmoid_table_205_3_sva_dfm_1;
  wire sigmoid_table_206_3_sva_dfm_1;
  wire sigmoid_table_207_3_sva_dfm_1;
  wire sigmoid_table_208_3_sva_dfm_1;
  wire sigmoid_table_209_3_sva_dfm_1;
  wire sigmoid_table_210_3_sva_dfm_1;
  wire sigmoid_table_211_3_sva_dfm_1;
  wire sigmoid_table_212_3_sva_dfm_1;
  wire sigmoid_table_213_3_sva_dfm_1;
  wire sigmoid_table_214_3_sva_dfm_1;
  wire sigmoid_table_215_3_sva_dfm_1;
  wire sigmoid_table_216_3_sva_dfm_1;
  wire sigmoid_table_217_3_sva_dfm_1;
  wire sigmoid_table_218_3_sva_dfm_1;
  wire sigmoid_table_219_3_sva_dfm_1;
  wire sigmoid_table_220_3_sva_dfm_1;
  wire sigmoid_table_221_3_sva_dfm_1;
  wire sigmoid_table_222_3_sva_dfm_1;
  wire sigmoid_table_223_3_sva_dfm_1;
  wire sigmoid_table_224_3_sva_dfm_1;
  wire sigmoid_table_225_3_sva_dfm_1;
  wire sigmoid_table_226_3_sva_dfm_1;
  wire sigmoid_table_227_3_sva_dfm_1;
  wire sigmoid_table_228_3_sva_dfm_1;
  wire sigmoid_table_274_3_sva_dfm_1;
  wire sigmoid_table_275_3_sva_dfm_1;
  wire sigmoid_table_276_3_sva_dfm_1;
  wire sigmoid_table_277_3_sva_dfm_1;
  wire sigmoid_table_278_3_sva_dfm_1;
  wire sigmoid_table_279_3_sva_dfm_1;
  wire sigmoid_table_280_3_sva_dfm_1;
  wire sigmoid_table_281_3_sva_dfm_1;
  wire sigmoid_table_282_3_sva_dfm_1;
  wire sigmoid_table_283_3_sva_dfm_1;
  wire sigmoid_table_308_3_sva_dfm_1;
  wire sigmoid_table_309_3_sva_dfm_1;
  wire sigmoid_table_310_3_sva_dfm_1;
  wire sigmoid_table_311_3_sva_dfm_1;
  wire sigmoid_table_312_3_sva_dfm_1;
  wire sigmoid_table_313_3_sva_dfm_1;
  wire sigmoid_table_330_3_sva_dfm_1;
  wire sigmoid_table_331_3_sva_dfm_1;
  wire sigmoid_table_332_3_sva_dfm_1;
  wire sigmoid_table_333_3_sva_dfm_1;
  wire sigmoid_table_334_3_sva_dfm_1;
  wire sigmoid_table_347_3_sva_dfm_1;
  wire sigmoid_table_348_3_sva_dfm_1;
  wire sigmoid_table_349_3_sva_dfm_1;
  wire sigmoid_table_350_3_sva_dfm_1;
  wire sigmoid_table_361_3_sva_dfm_1;
  wire sigmoid_table_362_3_sva_dfm_1;
  wire sigmoid_table_363_3_sva_dfm_1;
  wire sigmoid_table_373_3_sva_dfm_1;
  wire sigmoid_table_374_3_sva_dfm_1;
  wire sigmoid_table_375_3_sva_dfm_1;
  wire sigmoid_table_383_3_sva_dfm_1;
  wire sigmoid_table_384_3_sva_dfm_1;
  wire sigmoid_table_385_3_sva_dfm_1;
  wire sigmoid_table_392_3_sva_dfm_1;
  wire sigmoid_table_393_3_sva_dfm_1;
  wire sigmoid_table_394_3_sva_dfm_1;
  wire sigmoid_table_401_3_sva_dfm_1;
  wire sigmoid_table_402_3_sva_dfm_1;
  wire sigmoid_table_408_3_sva_dfm_1;
  wire sigmoid_table_409_3_sva_dfm_1;
  wire sigmoid_table_415_3_sva_dfm_1;
  wire sigmoid_table_416_3_sva_dfm_1;
  wire sigmoid_table_422_3_sva_dfm_1;
  wire sigmoid_table_428_3_sva_dfm_1;
  wire sigmoid_table_429_3_sva_dfm_1;
  wire sigmoid_table_434_3_sva_dfm_1;
  wire sigmoid_table_445_3_sva_dfm_1;
  wire sigmoid_table_450_3_sva_dfm_1;
  wire sigmoid_table_455_3_sva_dfm_1;
  wire sigmoid_table_460_3_sva_dfm_1;
  wire sigmoid_table_464_3_sva_dfm_1;
  wire sigmoid_table_469_3_sva_dfm_1;
  wire sigmoid_table_473_3_sva_dfm_1;
  wire sigmoid_table_478_3_sva_dfm_1;
  wire sigmoid_table_482_3_sva_dfm_1;
  wire sigmoid_table_486_3_sva_dfm_1;
  wire sigmoid_table_490_3_sva_dfm_1;
  wire sigmoid_table_494_3_sva_dfm_1;
  wire sigmoid_table_498_3_sva_dfm_1;
  wire sigmoid_table_502_3_sva_dfm_1;
  wire sigmoid_table_506_3_sva_dfm_1;
  wire sigmoid_table_514_3_sva_dfm_1;
  wire sigmoid_table_519_3_sva_dfm_1;
  wire sigmoid_table_523_3_sva_dfm_1;
  wire sigmoid_table_527_3_sva_dfm_1;
  wire sigmoid_table_531_3_sva_dfm_1;
  wire sigmoid_table_535_3_sva_dfm_1;
  wire sigmoid_table_539_3_sva_dfm_1;
  wire sigmoid_table_543_3_sva_dfm_1;
  wire sigmoid_table_547_3_sva_dfm_1;
  wire sigmoid_table_552_3_sva_dfm_1;
  wire sigmoid_table_556_3_sva_dfm_1;
  wire sigmoid_table_561_3_sva_dfm_1;
  wire sigmoid_table_565_3_sva_dfm_1;
  wire sigmoid_table_570_3_sva_dfm_1;
  wire sigmoid_table_575_3_sva_dfm_1;
  wire sigmoid_table_586_3_sva_dfm_1;
  wire sigmoid_table_591_3_sva_dfm_1;
  wire sigmoid_table_592_3_sva_dfm_1;
  wire sigmoid_table_597_3_sva_dfm_1;
  wire sigmoid_table_603_3_sva_dfm_1;
  wire sigmoid_table_604_3_sva_dfm_1;
  wire sigmoid_table_610_3_sva_dfm_1;
  wire sigmoid_table_617_3_sva_dfm_1;
  wire sigmoid_table_618_3_sva_dfm_1;
  wire sigmoid_table_624_3_sva_dfm_1;
  wire sigmoid_table_625_3_sva_dfm_1;
  wire sigmoid_table_633_3_sva_dfm_1;
  wire sigmoid_table_634_3_sva_dfm_1;
  wire sigmoid_table_642_3_sva_dfm_1;
  wire sigmoid_table_643_3_sva_dfm_1;
  wire sigmoid_table_652_3_sva_dfm_1;
  wire sigmoid_table_653_3_sva_dfm_1;
  wire sigmoid_table_654_3_sva_dfm_1;
  wire sigmoid_table_664_3_sva_dfm_1;
  wire sigmoid_table_665_3_sva_dfm_1;
  wire sigmoid_table_666_3_sva_dfm_1;
  wire sigmoid_table_678_3_sva_dfm_1;
  wire sigmoid_table_679_3_sva_dfm_1;
  wire sigmoid_table_680_3_sva_dfm_1;
  wire sigmoid_table_681_3_sva_dfm_1;
  wire sigmoid_table_695_3_sva_dfm_1;
  wire sigmoid_table_696_3_sva_dfm_1;
  wire sigmoid_table_697_3_sva_dfm_1;
  wire sigmoid_table_698_3_sva_dfm_1;
  wire sigmoid_table_699_3_sva_dfm_1;
  wire sigmoid_table_717_3_sva_dfm_1;
  wire sigmoid_table_718_3_sva_dfm_1;
  wire sigmoid_table_719_3_sva_dfm_1;
  wire sigmoid_table_720_3_sva_dfm_1;
  wire sigmoid_table_721_3_sva_dfm_1;
  wire sigmoid_table_722_3_sva_dfm_1;
  wire sigmoid_table_723_3_sva_dfm_1;
  wire sigmoid_table_751_3_sva_dfm_1;
  wire sigmoid_table_752_3_sva_dfm_1;
  wire sigmoid_table_753_3_sva_dfm_1;
  wire sigmoid_table_754_3_sva_dfm_1;
  wire sigmoid_table_755_3_sva_dfm_1;
  wire sigmoid_table_756_3_sva_dfm_1;
  wire sigmoid_table_757_3_sva_dfm_1;
  wire sigmoid_table_758_3_sva_dfm_1;
  wire sigmoid_table_759_3_sva_dfm_1;
  wire sigmoid_table_760_3_sva_dfm_1;
  wire sigmoid_table_761_3_sva_dfm_1;
  wire sigmoid_table_762_3_sva_dfm_1;
  wire sigmoid_table_339_6_sva_dfm_1;
  wire sigmoid_table_340_6_sva_dfm_1;
  wire sigmoid_table_341_6_sva_dfm_1;
  wire sigmoid_table_342_6_sva_dfm_1;
  wire sigmoid_table_343_6_sva_dfm_1;
  wire sigmoid_table_344_6_sva_dfm_1;
  wire sigmoid_table_345_6_sva_dfm_1;
  wire sigmoid_table_346_6_sva_dfm_1;
  wire sigmoid_table_347_6_sva_dfm_1;
  wire sigmoid_table_348_6_sva_dfm_1;
  wire sigmoid_table_349_6_sva_dfm_1;
  wire sigmoid_table_350_6_sva_dfm_1;
  wire sigmoid_table_351_6_sva_dfm_1;
  wire sigmoid_table_352_6_sva_dfm_1;
  wire sigmoid_table_353_6_sva_dfm_1;
  wire sigmoid_table_354_6_sva_dfm_1;
  wire sigmoid_table_355_6_sva_dfm_1;
  wire sigmoid_table_356_6_sva_dfm_1;
  wire sigmoid_table_357_6_sva_dfm_1;
  wire sigmoid_table_358_6_sva_dfm_1;
  wire sigmoid_table_359_6_sva_dfm_1;
  wire sigmoid_table_360_6_sva_dfm_1;
  wire sigmoid_table_361_6_sva_dfm_1;
  wire sigmoid_table_362_6_sva_dfm_1;
  wire sigmoid_table_363_6_sva_dfm_1;
  wire sigmoid_table_364_6_sva_dfm_1;
  wire sigmoid_table_365_6_sva_dfm_1;
  wire sigmoid_table_366_6_sva_dfm_1;
  wire sigmoid_table_367_5_sva_dfm_1;
  wire sigmoid_table_368_5_sva_dfm_1;
  wire sigmoid_table_369_5_sva_dfm_1;
  wire sigmoid_table_370_5_sva_dfm_1;
  wire sigmoid_table_371_5_sva_dfm_1;
  wire sigmoid_table_372_5_sva_dfm_1;
  wire sigmoid_table_373_5_sva_dfm_1;
  wire sigmoid_table_374_5_sva_dfm_1;
  wire sigmoid_table_375_5_sva_dfm_1;
  wire sigmoid_table_376_5_sva_dfm_1;
  wire sigmoid_table_377_5_sva_dfm_1;
  wire sigmoid_table_378_4_sva_dfm_1;
  wire sigmoid_table_379_4_sva_dfm_1;
  wire sigmoid_table_380_4_sva_dfm_1;
  wire sigmoid_table_381_4_sva_dfm_1;
  wire sigmoid_table_382_4_sva_dfm_1;
  wire sigmoid_table_462_6_sva_dfm_1;
  wire sigmoid_table_463_6_sva_dfm_1;
  wire sigmoid_table_464_6_sva_dfm_1;
  wire sigmoid_table_465_6_sva_dfm_1;
  wire sigmoid_table_466_6_sva_dfm_1;
  wire sigmoid_table_467_6_sva_dfm_1;
  wire sigmoid_table_468_6_sva_dfm_1;
  wire sigmoid_table_469_6_sva_dfm_1;
  wire sigmoid_table_470_6_sva_dfm_1;
  wire sigmoid_table_471_5_sva_dfm_1;
  wire sigmoid_table_472_5_sva_dfm_1;
  wire sigmoid_table_473_5_sva_dfm_1;
  wire sigmoid_table_474_5_sva_dfm_1;
  wire sigmoid_table_475_5_sva_dfm_1;
  wire sigmoid_table_476_4_sva_dfm_1;
  wire sigmoid_table_477_4_sva_dfm_1;
  wire sigmoid_table_529_6_sva_dfm_1;
  wire sigmoid_table_530_6_sva_dfm_1;
  wire sigmoid_table_531_6_sva_dfm_1;
  wire sigmoid_table_532_6_sva_dfm_1;
  wire sigmoid_table_533_6_sva_dfm_1;
  wire sigmoid_table_534_6_sva_dfm_1;
  wire sigmoid_table_535_6_sva_dfm_1;
  wire sigmoid_table_536_6_sva_dfm_1;
  wire sigmoid_table_537_5_sva_dfm_1;
  wire sigmoid_table_538_5_sva_dfm_1;
  wire sigmoid_table_539_5_sva_dfm_1;
  wire sigmoid_table_540_5_sva_dfm_1;
  wire sigmoid_table_541_4_sva_dfm_1;
  wire sigmoid_table_542_4_sva_dfm_1;
  wire sigmoid_table_606_6_sva_dfm_1;
  wire sigmoid_table_607_6_sva_dfm_1;
  wire sigmoid_table_608_6_sva_dfm_1;
  wire sigmoid_table_609_6_sva_dfm_1;
  wire sigmoid_table_610_6_sva_dfm_1;
  wire sigmoid_table_611_6_sva_dfm_1;
  wire sigmoid_table_612_6_sva_dfm_1;
  wire sigmoid_table_613_6_sva_dfm_1;
  wire sigmoid_table_614_6_sva_dfm_1;
  wire sigmoid_table_615_6_sva_dfm_1;
  wire sigmoid_table_616_6_sva_dfm_1;
  wire sigmoid_table_617_6_sva_dfm_1;
  wire sigmoid_table_618_6_sva_dfm_1;
  wire sigmoid_table_619_6_sva_dfm_1;
  wire sigmoid_table_620_5_sva_dfm_1;
  wire sigmoid_table_621_5_sva_dfm_1;
  wire sigmoid_table_622_5_sva_dfm_1;
  wire sigmoid_table_623_5_sva_dfm_1;
  wire sigmoid_table_624_5_sva_dfm_1;
  wire sigmoid_table_625_5_sva_dfm_1;
  wire sigmoid_table_626_5_sva_dfm_1;
  wire sigmoid_table_627_5_sva_dfm_1;
  wire sigmoid_table_628_4_sva_dfm_1;
  wire sigmoid_table_629_4_sva_dfm_1;
  wire sigmoid_table_630_4_sva_dfm_1;
  wire sigmoid_table_631_4_sva_dfm_1;
  wire sigmoid_table_632_4_sva_dfm_1;
  wire sigmoid_table_247_4_sva_dfm_1;
  wire sigmoid_table_248_4_sva_dfm_1;
  wire sigmoid_table_249_4_sva_dfm_1;
  wire sigmoid_table_250_4_sva_dfm_1;
  wire sigmoid_table_251_4_sva_dfm_1;
  wire sigmoid_table_252_4_sva_dfm_1;
  wire sigmoid_table_253_4_sva_dfm_1;
  wire sigmoid_table_254_4_sva_dfm_1;
  wire sigmoid_table_255_4_sva_dfm_1;
  wire sigmoid_table_256_4_sva_dfm_1;
  wire sigmoid_table_257_4_sva_dfm_1;
  wire sigmoid_table_258_4_sva_dfm_1;
  wire sigmoid_table_259_4_sva_dfm_1;
  wire sigmoid_table_260_4_sva_dfm_1;
  wire sigmoid_table_261_4_sva_dfm_1;
  wire sigmoid_table_262_4_sva_dfm_1;
  wire sigmoid_table_263_4_sva_dfm_1;
  wire sigmoid_table_264_4_sva_dfm_1;
  wire sigmoid_table_265_4_sva_dfm_1;
  wire sigmoid_table_266_4_sva_dfm_1;
  wire sigmoid_table_267_4_sva_dfm_1;
  wire sigmoid_table_268_4_sva_dfm_1;
  wire sigmoid_table_269_4_sva_dfm_1;
  wire sigmoid_table_270_4_sva_dfm_1;
  wire sigmoid_table_271_4_sva_dfm_1;
  wire sigmoid_table_272_4_sva_dfm_1;
  wire sigmoid_table_273_4_sva_dfm_1;
  wire sigmoid_table_320_4_sva_dfm_1;
  wire sigmoid_table_321_4_sva_dfm_1;
  wire sigmoid_table_322_4_sva_dfm_1;
  wire sigmoid_table_323_4_sva_dfm_1;
  wire sigmoid_table_324_4_sva_dfm_1;
  wire sigmoid_table_325_4_sva_dfm_1;
  wire sigmoid_table_326_4_sva_dfm_1;
  wire sigmoid_table_327_4_sva_dfm_1;
  wire sigmoid_table_328_4_sva_dfm_1;
  wire sigmoid_table_329_4_sva_dfm_1;
  wire sigmoid_table_355_4_sva_dfm_1;
  wire sigmoid_table_356_4_sva_dfm_1;
  wire sigmoid_table_357_4_sva_dfm_1;
  wire sigmoid_table_358_4_sva_dfm_1;
  wire sigmoid_table_359_4_sva_dfm_1;
  wire sigmoid_table_360_4_sva_dfm_1;
  wire sigmoid_table_397_4_sva_dfm_1;
  wire sigmoid_table_398_4_sva_dfm_1;
  wire sigmoid_table_399_4_sva_dfm_1;
  wire sigmoid_table_400_4_sva_dfm_1;
  wire sigmoid_table_412_4_sva_dfm_1;
  wire sigmoid_table_413_4_sva_dfm_1;
  wire sigmoid_table_414_4_sva_dfm_1;
  wire sigmoid_table_425_4_sva_dfm_1;
  wire sigmoid_table_426_4_sva_dfm_1;
  wire sigmoid_table_427_4_sva_dfm_1;
  wire sigmoid_table_447_4_sva_dfm_1;
  wire sigmoid_table_448_4_sva_dfm_1;
  wire sigmoid_table_449_4_sva_dfm_1;
  wire sigmoid_table_457_4_sva_dfm_1;
  wire sigmoid_table_458_4_sva_dfm_1;
  wire sigmoid_table_459_4_sva_dfm_1;
  wire sigmoid_table_467_4_sva_dfm_1;
  wire sigmoid_table_468_4_sva_dfm_1;
  wire sigmoid_table_484_4_sva_dfm_1;
  wire sigmoid_table_485_4_sva_dfm_1;
  wire sigmoid_table_492_4_sva_dfm_1;
  wire sigmoid_table_493_4_sva_dfm_1;
  wire sigmoid_table_500_4_sva_dfm_1;
  wire sigmoid_table_501_4_sva_dfm_1;
  wire sigmoid_table_517_4_sva_dfm_1;
  wire sigmoid_table_518_4_sva_dfm_1;
  wire sigmoid_table_525_4_sva_dfm_1;
  wire sigmoid_table_526_4_sva_dfm_1;
  wire sigmoid_table_533_4_sva_dfm_1;
  wire sigmoid_table_534_4_sva_dfm_1;
  wire sigmoid_table_549_4_sva_dfm_1;
  wire sigmoid_table_550_4_sva_dfm_1;
  wire sigmoid_table_551_4_sva_dfm_1;
  wire sigmoid_table_558_4_sva_dfm_1;
  wire sigmoid_table_559_4_sva_dfm_1;
  wire sigmoid_table_560_4_sva_dfm_1;
  wire sigmoid_table_568_4_sva_dfm_1;
  wire sigmoid_table_569_4_sva_dfm_1;
  wire sigmoid_table_588_4_sva_dfm_1;
  wire sigmoid_table_589_4_sva_dfm_1;
  wire sigmoid_table_590_4_sva_dfm_1;
  wire sigmoid_table_600_4_sva_dfm_1;
  wire sigmoid_table_601_4_sva_dfm_1;
  wire sigmoid_table_602_4_sva_dfm_1;
  wire sigmoid_table_613_4_sva_dfm_1;
  wire sigmoid_table_614_4_sva_dfm_1;
  wire sigmoid_table_615_4_sva_dfm_1;
  wire sigmoid_table_616_4_sva_dfm_1;
  wire sigmoid_table_647_4_sva_dfm_1;
  wire sigmoid_table_648_4_sva_dfm_1;
  wire sigmoid_table_649_4_sva_dfm_1;
  wire sigmoid_table_650_4_sva_dfm_1;
  wire sigmoid_table_651_4_sva_dfm_1;
  wire sigmoid_table_670_4_sva_dfm_1;
  wire sigmoid_table_671_4_sva_dfm_1;
  wire sigmoid_table_672_4_sva_dfm_1;
  wire sigmoid_table_673_4_sva_dfm_1;
  wire sigmoid_table_674_4_sva_dfm_1;
  wire sigmoid_table_675_4_sva_dfm_1;
  wire sigmoid_table_676_4_sva_dfm_1;
  wire sigmoid_table_677_4_sva_dfm_1;
  wire sigmoid_table_705_4_sva_dfm_1;
  wire sigmoid_table_706_4_sva_dfm_1;
  wire sigmoid_table_707_4_sva_dfm_1;
  wire sigmoid_table_708_4_sva_dfm_1;
  wire sigmoid_table_709_4_sva_dfm_1;
  wire sigmoid_table_710_4_sva_dfm_1;
  wire sigmoid_table_711_4_sva_dfm_1;
  wire sigmoid_table_712_4_sva_dfm_1;
  wire sigmoid_table_713_4_sva_dfm_1;
  wire sigmoid_table_714_4_sva_dfm_1;
  wire sigmoid_table_715_4_sva_dfm_1;
  wire sigmoid_table_716_4_sva_dfm_1;
  wire sigmoid_table_293_5_sva_dfm_1;
  wire sigmoid_table_294_5_sva_dfm_1;
  wire sigmoid_table_295_5_sva_dfm_1;
  wire sigmoid_table_296_5_sva_dfm_1;
  wire sigmoid_table_297_5_sva_dfm_1;
  wire sigmoid_table_298_5_sva_dfm_1;
  wire sigmoid_table_299_5_sva_dfm_1;
  wire sigmoid_table_300_5_sva_dfm_1;
  wire sigmoid_table_301_5_sva_dfm_1;
  wire sigmoid_table_302_5_sva_dfm_1;
  wire sigmoid_table_303_5_sva_dfm_1;
  wire sigmoid_table_304_5_sva_dfm_1;
  wire sigmoid_table_305_5_sva_dfm_1;
  wire sigmoid_table_306_5_sva_dfm_1;
  wire sigmoid_table_307_5_sva_dfm_1;
  wire sigmoid_table_308_5_sva_dfm_1;
  wire sigmoid_table_309_5_sva_dfm_1;
  wire sigmoid_table_310_5_sva_dfm_1;
  wire sigmoid_table_311_5_sva_dfm_1;
  wire sigmoid_table_312_5_sva_dfm_1;
  wire sigmoid_table_313_5_sva_dfm_1;
  wire sigmoid_table_314_5_sva_dfm_1;
  wire sigmoid_table_315_5_sva_dfm_1;
  wire sigmoid_table_316_5_sva_dfm_1;
  wire sigmoid_table_317_5_sva_dfm_1;
  wire sigmoid_table_318_5_sva_dfm_1;
  wire sigmoid_table_319_5_sva_dfm_1;
  wire sigmoid_table_405_5_sva_dfm_1;
  wire sigmoid_table_406_5_sva_dfm_1;
  wire sigmoid_table_407_5_sva_dfm_1;
  wire sigmoid_table_408_5_sva_dfm_1;
  wire sigmoid_table_409_5_sva_dfm_1;
  wire sigmoid_table_410_5_sva_dfm_1;
  wire sigmoid_table_411_5_sva_dfm_1;
  wire sigmoid_table_452_5_sva_dfm_1;
  wire sigmoid_table_453_5_sva_dfm_1;
  wire sigmoid_table_454_5_sva_dfm_1;
  wire sigmoid_table_455_5_sva_dfm_1;
  wire sigmoid_table_456_5_sva_dfm_1;
  wire sigmoid_table_488_5_sva_dfm_1;
  wire sigmoid_table_489_5_sva_dfm_1;
  wire sigmoid_table_490_5_sva_dfm_1;
  wire sigmoid_table_491_5_sva_dfm_1;
  wire sigmoid_table_521_5_sva_dfm_1;
  wire sigmoid_table_522_5_sva_dfm_1;
  wire sigmoid_table_523_5_sva_dfm_1;
  wire sigmoid_table_524_5_sva_dfm_1;
  wire sigmoid_table_554_5_sva_dfm_1;
  wire sigmoid_table_555_5_sva_dfm_1;
  wire sigmoid_table_556_5_sva_dfm_1;
  wire sigmoid_table_557_5_sva_dfm_1;
  wire sigmoid_table_594_5_sva_dfm_1;
  wire sigmoid_table_595_5_sva_dfm_1;
  wire sigmoid_table_596_5_sva_dfm_1;
  wire sigmoid_table_597_5_sva_dfm_1;
  wire sigmoid_table_598_5_sva_dfm_1;
  wire sigmoid_table_599_5_sva_dfm_1;
  wire sigmoid_table_658_5_sva_dfm_1;
  wire sigmoid_table_659_5_sva_dfm_1;
  wire sigmoid_table_660_5_sva_dfm_1;
  wire sigmoid_table_661_5_sva_dfm_1;
  wire sigmoid_table_662_5_sva_dfm_1;
  wire sigmoid_table_663_5_sva_dfm_1;
  wire sigmoid_table_664_5_sva_dfm_1;
  wire sigmoid_table_665_5_sva_dfm_1;
  wire sigmoid_table_666_5_sva_dfm_1;
  wire sigmoid_table_667_5_sva_dfm_1;
  wire sigmoid_table_668_5_sva_dfm_1;
  wire sigmoid_table_669_5_sva_dfm_1;
  wire [5:0] operator_32_true_acc_psp_sva_1;
  wire [6:0] nl_operator_32_true_acc_psp_sva_1;
  wire for_for_or_1_itm;
  wire [8:0] for_for_or_itm;
  wire operator_32_true_acc_itm_4;

  wire[4:0] operator_32_true_acc_nl;
  wire[5:0] nl_operator_32_true_acc_nl;
  wire[0:0] operator_32_true_not_2_nl;
  wire[8:0] for_for_and_1_nl;
  wire[0:0] operator_32_true_not_4_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [17:0] nl_res_rsci_d;
  assign nl_res_rsci_d = {8'b00000000 , res_rsci_d_9 , res_rsci_d_8 , res_rsci_d_7
      , res_rsci_d_6 , res_rsci_d_5 , res_rsci_d_4 , res_rsci_d_3 , res_rsci_d_2
      , res_rsci_d_1 , res_rsci_d_0};
  ccs_in_v1 #(.rscid(32'sd13),
  .width(32'sd18)) data_rsci (
      .dat(data_rsc_dat),
      .idat(data_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd14),
  .width(32'sd18)) res_rsci (
      .d(nl_res_rsci_d[17:0]),
      .z(res_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd27),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign sigmoid_table_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  assign sigmoid_table_69_0_sva_dfm_1 = sigmoid_table_69_0_sva | (~ initialized_sva);
  assign sigmoid_table_70_0_sva_dfm_1 = sigmoid_table_70_0_sva | (~ initialized_sva);
  assign sigmoid_table_71_0_sva_dfm_1 = sigmoid_table_71_0_sva | (~ initialized_sva);
  assign sigmoid_table_72_0_sva_dfm_1 = sigmoid_table_72_0_sva | (~ initialized_sva);
  assign sigmoid_table_73_0_sva_dfm_1 = sigmoid_table_73_0_sva | (~ initialized_sva);
  assign sigmoid_table_74_0_sva_dfm_1 = sigmoid_table_74_0_sva | (~ initialized_sva);
  assign sigmoid_table_75_0_sva_dfm_1 = sigmoid_table_75_0_sva | (~ initialized_sva);
  assign sigmoid_table_76_0_sva_dfm_1 = sigmoid_table_76_0_sva | (~ initialized_sva);
  assign sigmoid_table_77_0_sva_dfm_1 = sigmoid_table_77_0_sva | (~ initialized_sva);
  assign sigmoid_table_78_0_sva_dfm_1 = sigmoid_table_78_0_sva | (~ initialized_sva);
  assign sigmoid_table_79_0_sva_dfm_1 = sigmoid_table_79_0_sva | (~ initialized_sva);
  assign sigmoid_table_80_0_sva_dfm_1 = sigmoid_table_80_0_sva | (~ initialized_sva);
  assign sigmoid_table_81_0_sva_dfm_1 = sigmoid_table_81_0_sva | (~ initialized_sva);
  assign sigmoid_table_82_0_sva_dfm_1 = sigmoid_table_82_0_sva | (~ initialized_sva);
  assign sigmoid_table_83_0_sva_dfm_1 = sigmoid_table_83_0_sva | (~ initialized_sva);
  assign sigmoid_table_84_0_sva_dfm_1 = sigmoid_table_84_0_sva | (~ initialized_sva);
  assign sigmoid_table_85_0_sva_dfm_1 = sigmoid_table_85_0_sva | (~ initialized_sva);
  assign sigmoid_table_86_0_sva_dfm_1 = sigmoid_table_86_0_sva | (~ initialized_sva);
  assign sigmoid_table_87_0_sva_dfm_1 = sigmoid_table_87_0_sva | (~ initialized_sva);
  assign sigmoid_table_88_0_sva_dfm_1 = sigmoid_table_88_0_sva | (~ initialized_sva);
  assign sigmoid_table_89_0_sva_dfm_1 = sigmoid_table_89_0_sva | (~ initialized_sva);
  assign sigmoid_table_90_0_sva_dfm_1 = sigmoid_table_90_0_sva | (~ initialized_sva);
  assign sigmoid_table_91_0_sva_dfm_1 = sigmoid_table_91_0_sva | (~ initialized_sva);
  assign sigmoid_table_92_0_sva_dfm_1 = sigmoid_table_92_0_sva | (~ initialized_sva);
  assign sigmoid_table_93_0_sva_dfm_1 = sigmoid_table_93_0_sva | (~ initialized_sva);
  assign sigmoid_table_94_0_sva_dfm_1 = sigmoid_table_94_0_sva | (~ initialized_sva);
  assign sigmoid_table_95_0_sva_dfm_1 = sigmoid_table_95_0_sva | (~ initialized_sva);
  assign sigmoid_table_96_0_sva_dfm_1 = sigmoid_table_96_0_sva | (~ initialized_sva);
  assign sigmoid_table_97_0_sva_dfm_1 = sigmoid_table_97_0_sva | (~ initialized_sva);
  assign sigmoid_table_98_0_sva_dfm_1 = sigmoid_table_98_0_sva | (~ initialized_sva);
  assign sigmoid_table_99_0_sva_dfm_1 = sigmoid_table_99_0_sva | (~ initialized_sva);
  assign sigmoid_table_100_0_sva_dfm_1 = sigmoid_table_100_0_sva | (~ initialized_sva);
  assign sigmoid_table_101_0_sva_dfm_1 = sigmoid_table_101_0_sva | (~ initialized_sva);
  assign sigmoid_table_102_0_sva_dfm_1 = sigmoid_table_102_0_sva | (~ initialized_sva);
  assign sigmoid_table_103_0_sva_dfm_1 = sigmoid_table_103_0_sva | (~ initialized_sva);
  assign sigmoid_table_104_0_sva_dfm_1 = sigmoid_table_104_0_sva | (~ initialized_sva);
  assign sigmoid_table_105_0_sva_dfm_1 = sigmoid_table_105_0_sva | (~ initialized_sva);
  assign sigmoid_table_106_0_sva_dfm_1 = sigmoid_table_106_0_sva | (~ initialized_sva);
  assign sigmoid_table_107_0_sva_dfm_1 = sigmoid_table_107_0_sva | (~ initialized_sva);
  assign sigmoid_table_108_0_sva_dfm_1 = sigmoid_table_108_0_sva | (~ initialized_sva);
  assign sigmoid_table_109_0_sva_dfm_1 = sigmoid_table_109_0_sva | (~ initialized_sva);
  assign sigmoid_table_110_0_sva_dfm_1 = sigmoid_table_110_0_sva | (~ initialized_sva);
  assign sigmoid_table_111_0_sva_dfm_1 = sigmoid_table_111_0_sva | (~ initialized_sva);
  assign sigmoid_table_112_0_sva_dfm_1 = sigmoid_table_112_0_sva | (~ initialized_sva);
  assign sigmoid_table_139_0_sva_dfm_1 = sigmoid_table_139_0_sva | (~ initialized_sva);
  assign sigmoid_table_140_0_sva_dfm_1 = sigmoid_table_140_0_sva | (~ initialized_sva);
  assign sigmoid_table_141_0_sva_dfm_1 = sigmoid_table_141_0_sva | (~ initialized_sva);
  assign sigmoid_table_142_0_sva_dfm_1 = sigmoid_table_142_0_sva | (~ initialized_sva);
  assign sigmoid_table_143_0_sva_dfm_1 = sigmoid_table_143_0_sva | (~ initialized_sva);
  assign sigmoid_table_144_0_sva_dfm_1 = sigmoid_table_144_0_sva | (~ initialized_sva);
  assign sigmoid_table_145_0_sva_dfm_1 = sigmoid_table_145_0_sva | (~ initialized_sva);
  assign sigmoid_table_146_0_sva_dfm_1 = sigmoid_table_146_0_sva | (~ initialized_sva);
  assign sigmoid_table_147_0_sva_dfm_1 = sigmoid_table_147_0_sva | (~ initialized_sva);
  assign sigmoid_table_148_0_sva_dfm_1 = sigmoid_table_148_0_sva | (~ initialized_sva);
  assign sigmoid_table_149_0_sva_dfm_1 = sigmoid_table_149_0_sva | (~ initialized_sva);
  assign sigmoid_table_150_0_sva_dfm_1 = sigmoid_table_150_0_sva | (~ initialized_sva);
  assign sigmoid_table_151_0_sva_dfm_1 = sigmoid_table_151_0_sva | (~ initialized_sva);
  assign sigmoid_table_152_0_sva_dfm_1 = sigmoid_table_152_0_sva | (~ initialized_sva);
  assign sigmoid_table_153_0_sva_dfm_1 = sigmoid_table_153_0_sva | (~ initialized_sva);
  assign sigmoid_table_154_0_sva_dfm_1 = sigmoid_table_154_0_sva | (~ initialized_sva);
  assign sigmoid_table_155_0_sva_dfm_1 = sigmoid_table_155_0_sva | (~ initialized_sva);
  assign sigmoid_table_156_0_sva_dfm_1 = sigmoid_table_156_0_sva | (~ initialized_sva);
  assign sigmoid_table_157_0_sva_dfm_1 = sigmoid_table_157_0_sva | (~ initialized_sva);
  assign sigmoid_table_172_0_sva_dfm_1 = sigmoid_table_172_0_sva | (~ initialized_sva);
  assign sigmoid_table_173_0_sva_dfm_1 = sigmoid_table_173_0_sva | (~ initialized_sva);
  assign sigmoid_table_174_0_sva_dfm_1 = sigmoid_table_174_0_sva | (~ initialized_sva);
  assign sigmoid_table_175_0_sva_dfm_1 = sigmoid_table_175_0_sva | (~ initialized_sva);
  assign sigmoid_table_176_0_sva_dfm_1 = sigmoid_table_176_0_sva | (~ initialized_sva);
  assign sigmoid_table_177_0_sva_dfm_1 = sigmoid_table_177_0_sva | (~ initialized_sva);
  assign sigmoid_table_178_0_sva_dfm_1 = sigmoid_table_178_0_sva | (~ initialized_sva);
  assign sigmoid_table_179_0_sva_dfm_1 = sigmoid_table_179_0_sva | (~ initialized_sva);
  assign sigmoid_table_180_0_sva_dfm_1 = sigmoid_table_180_0_sva | (~ initialized_sva);
  assign sigmoid_table_181_0_sva_dfm_1 = sigmoid_table_181_0_sva | (~ initialized_sva);
  assign sigmoid_table_182_0_sva_dfm_1 = sigmoid_table_182_0_sva | (~ initialized_sva);
  assign sigmoid_table_183_0_sva_dfm_1 = sigmoid_table_183_0_sva | (~ initialized_sva);
  assign sigmoid_table_194_0_sva_dfm_1 = sigmoid_table_194_0_sva | (~ initialized_sva);
  assign sigmoid_table_195_0_sva_dfm_1 = sigmoid_table_195_0_sva | (~ initialized_sva);
  assign sigmoid_table_196_0_sva_dfm_1 = sigmoid_table_196_0_sva | (~ initialized_sva);
  assign sigmoid_table_197_0_sva_dfm_1 = sigmoid_table_197_0_sva | (~ initialized_sva);
  assign sigmoid_table_198_0_sva_dfm_1 = sigmoid_table_198_0_sva | (~ initialized_sva);
  assign sigmoid_table_199_0_sva_dfm_1 = sigmoid_table_199_0_sva | (~ initialized_sva);
  assign sigmoid_table_200_0_sva_dfm_1 = sigmoid_table_200_0_sva | (~ initialized_sva);
  assign sigmoid_table_201_0_sva_dfm_1 = sigmoid_table_201_0_sva | (~ initialized_sva);
  assign sigmoid_table_210_0_sva_dfm_1 = sigmoid_table_210_0_sva | (~ initialized_sva);
  assign sigmoid_table_211_0_sva_dfm_1 = sigmoid_table_211_0_sva | (~ initialized_sva);
  assign sigmoid_table_212_0_sva_dfm_1 = sigmoid_table_212_0_sva | (~ initialized_sva);
  assign sigmoid_table_213_0_sva_dfm_1 = sigmoid_table_213_0_sva | (~ initialized_sva);
  assign sigmoid_table_214_0_sva_dfm_1 = sigmoid_table_214_0_sva | (~ initialized_sva);
  assign sigmoid_table_215_0_sva_dfm_1 = sigmoid_table_215_0_sva | (~ initialized_sva);
  assign sigmoid_table_216_0_sva_dfm_1 = sigmoid_table_216_0_sva | (~ initialized_sva);
  assign sigmoid_table_223_0_sva_dfm_1 = sigmoid_table_223_0_sva | (~ initialized_sva);
  assign sigmoid_table_224_0_sva_dfm_1 = sigmoid_table_224_0_sva | (~ initialized_sva);
  assign sigmoid_table_225_0_sva_dfm_1 = sigmoid_table_225_0_sva | (~ initialized_sva);
  assign sigmoid_table_226_0_sva_dfm_1 = sigmoid_table_226_0_sva | (~ initialized_sva);
  assign sigmoid_table_227_0_sva_dfm_1 = sigmoid_table_227_0_sva | (~ initialized_sva);
  assign sigmoid_table_228_0_sva_dfm_1 = sigmoid_table_228_0_sva | (~ initialized_sva);
  assign sigmoid_table_234_0_sva_dfm_1 = sigmoid_table_234_0_sva | (~ initialized_sva);
  assign sigmoid_table_235_0_sva_dfm_1 = sigmoid_table_235_0_sva | (~ initialized_sva);
  assign sigmoid_table_236_0_sva_dfm_1 = sigmoid_table_236_0_sva | (~ initialized_sva);
  assign sigmoid_table_237_0_sva_dfm_1 = sigmoid_table_237_0_sva | (~ initialized_sva);
  assign sigmoid_table_238_0_sva_dfm_1 = sigmoid_table_238_0_sva | (~ initialized_sva);
  assign sigmoid_table_243_0_sva_dfm_1 = sigmoid_table_243_0_sva | (~ initialized_sva);
  assign sigmoid_table_244_0_sva_dfm_1 = sigmoid_table_244_0_sva | (~ initialized_sva);
  assign sigmoid_table_245_0_sva_dfm_1 = sigmoid_table_245_0_sva | (~ initialized_sva);
  assign sigmoid_table_246_0_sva_dfm_1 = sigmoid_table_246_0_sva | (~ initialized_sva);
  assign sigmoid_table_251_0_sva_dfm_1 = sigmoid_table_251_0_sva | (~ initialized_sva);
  assign sigmoid_table_252_0_sva_dfm_1 = sigmoid_table_252_0_sva | (~ initialized_sva);
  assign sigmoid_table_253_0_sva_dfm_1 = sigmoid_table_253_0_sva | (~ initialized_sva);
  assign sigmoid_table_254_0_sva_dfm_1 = sigmoid_table_254_0_sva | (~ initialized_sva);
  assign sigmoid_table_259_0_sva_dfm_1 = sigmoid_table_259_0_sva | (~ initialized_sva);
  assign sigmoid_table_260_0_sva_dfm_1 = sigmoid_table_260_0_sva | (~ initialized_sva);
  assign sigmoid_table_261_0_sva_dfm_1 = sigmoid_table_261_0_sva | (~ initialized_sva);
  assign sigmoid_table_265_0_sva_dfm_1 = sigmoid_table_265_0_sva | (~ initialized_sva);
  assign sigmoid_table_266_0_sva_dfm_1 = sigmoid_table_266_0_sva | (~ initialized_sva);
  assign sigmoid_table_267_0_sva_dfm_1 = sigmoid_table_267_0_sva | (~ initialized_sva);
  assign sigmoid_table_271_0_sva_dfm_1 = sigmoid_table_271_0_sva | (~ initialized_sva);
  assign sigmoid_table_272_0_sva_dfm_1 = sigmoid_table_272_0_sva | (~ initialized_sva);
  assign sigmoid_table_273_0_sva_dfm_1 = sigmoid_table_273_0_sva | (~ initialized_sva);
  assign sigmoid_table_276_0_sva_dfm_1 = sigmoid_table_276_0_sva | (~ initialized_sva);
  assign sigmoid_table_277_0_sva_dfm_1 = sigmoid_table_277_0_sva | (~ initialized_sva);
  assign sigmoid_table_278_0_sva_dfm_1 = sigmoid_table_278_0_sva | (~ initialized_sva);
  assign sigmoid_table_282_0_sva_dfm_1 = sigmoid_table_282_0_sva | (~ initialized_sva);
  assign sigmoid_table_283_0_sva_dfm_1 = sigmoid_table_283_0_sva | (~ initialized_sva);
  assign sigmoid_table_286_0_sva_dfm_1 = sigmoid_table_286_0_sva | (~ initialized_sva);
  assign sigmoid_table_287_0_sva_dfm_1 = sigmoid_table_287_0_sva | (~ initialized_sva);
  assign sigmoid_table_291_0_sva_dfm_1 = sigmoid_table_291_0_sva | (~ initialized_sva);
  assign sigmoid_table_292_0_sva_dfm_1 = sigmoid_table_292_0_sva | (~ initialized_sva);
  assign sigmoid_table_295_0_sva_dfm_1 = sigmoid_table_295_0_sva | (~ initialized_sva);
  assign sigmoid_table_296_0_sva_dfm_1 = sigmoid_table_296_0_sva | (~ initialized_sva);
  assign sigmoid_table_299_0_sva_dfm_1 = sigmoid_table_299_0_sva | (~ initialized_sva);
  assign sigmoid_table_300_0_sva_dfm_1 = sigmoid_table_300_0_sva | (~ initialized_sva);
  assign sigmoid_table_302_0_sva_dfm_1 = sigmoid_table_302_0_sva | (~ initialized_sva);
  assign sigmoid_table_303_0_sva_dfm_1 = sigmoid_table_303_0_sva | (~ initialized_sva);
  assign sigmoid_table_306_0_sva_dfm_1 = sigmoid_table_306_0_sva | (~ initialized_sva);
  assign sigmoid_table_307_0_sva_dfm_1 = sigmoid_table_307_0_sva | (~ initialized_sva);
  assign sigmoid_table_309_0_sva_dfm_1 = sigmoid_table_309_0_sva | (~ initialized_sva);
  assign sigmoid_table_310_0_sva_dfm_1 = sigmoid_table_310_0_sva | (~ initialized_sva);
  assign sigmoid_table_312_0_sva_dfm_1 = sigmoid_table_312_0_sva | (~ initialized_sva);
  assign sigmoid_table_313_0_sva_dfm_1 = sigmoid_table_313_0_sva | (~ initialized_sva);
  assign sigmoid_table_315_0_sva_dfm_1 = sigmoid_table_315_0_sva | (~ initialized_sva);
  assign sigmoid_table_316_0_sva_dfm_1 = sigmoid_table_316_0_sva | (~ initialized_sva);
  assign sigmoid_table_318_0_sva_dfm_1 = sigmoid_table_318_0_sva | (~ initialized_sva);
  assign sigmoid_table_319_0_sva_dfm_1 = sigmoid_table_319_0_sva | (~ initialized_sva);
  assign sigmoid_table_321_0_sva_dfm_1 = sigmoid_table_321_0_sva | (~ initialized_sva);
  assign sigmoid_table_324_0_sva_dfm_1 = sigmoid_table_324_0_sva | (~ initialized_sva);
  assign sigmoid_table_326_0_sva_dfm_1 = sigmoid_table_326_0_sva | (~ initialized_sva);
  assign sigmoid_table_327_0_sva_dfm_1 = sigmoid_table_327_0_sva | (~ initialized_sva);
  assign sigmoid_table_329_0_sva_dfm_1 = sigmoid_table_329_0_sva | (~ initialized_sva);
  assign sigmoid_table_331_0_sva_dfm_1 = sigmoid_table_331_0_sva | (~ initialized_sva);
  assign sigmoid_table_334_0_sva_dfm_1 = sigmoid_table_334_0_sva | (~ initialized_sva);
  assign sigmoid_table_336_0_sva_dfm_1 = sigmoid_table_336_0_sva | (~ initialized_sva);
  assign sigmoid_table_338_0_sva_dfm_1 = sigmoid_table_338_0_sva | (~ initialized_sva);
  assign sigmoid_table_340_0_sva_dfm_1 = sigmoid_table_340_0_sva | (~ initialized_sva);
  assign sigmoid_table_342_0_sva_dfm_1 = sigmoid_table_342_0_sva | (~ initialized_sva);
  assign sigmoid_table_344_0_sva_dfm_1 = sigmoid_table_344_0_sva | (~ initialized_sva);
  assign sigmoid_table_346_0_sva_dfm_1 = sigmoid_table_346_0_sva | (~ initialized_sva);
  assign sigmoid_table_348_0_sva_dfm_1 = sigmoid_table_348_0_sva | (~ initialized_sva);
  assign sigmoid_table_350_0_sva_dfm_1 = sigmoid_table_350_0_sva | (~ initialized_sva);
  assign sigmoid_table_352_0_sva_dfm_1 = sigmoid_table_352_0_sva | (~ initialized_sva);
  assign sigmoid_table_354_0_sva_dfm_1 = sigmoid_table_354_0_sva | (~ initialized_sva);
  assign sigmoid_table_355_0_sva_dfm_1 = sigmoid_table_355_0_sva | (~ initialized_sva);
  assign sigmoid_table_357_0_sva_dfm_1 = sigmoid_table_357_0_sva | (~ initialized_sva);
  assign sigmoid_table_359_0_sva_dfm_1 = sigmoid_table_359_0_sva | (~ initialized_sva);
  assign sigmoid_table_360_0_sva_dfm_1 = sigmoid_table_360_0_sva | (~ initialized_sva);
  assign sigmoid_table_362_0_sva_dfm_1 = sigmoid_table_362_0_sva | (~ initialized_sva);
  assign sigmoid_table_365_0_sva_dfm_1 = sigmoid_table_365_0_sva | (~ initialized_sva);
  assign sigmoid_table_368_0_sva_dfm_1 = sigmoid_table_368_0_sva | (~ initialized_sva);
  assign sigmoid_table_369_0_sva_dfm_1 = sigmoid_table_369_0_sva | (~ initialized_sva);
  assign sigmoid_table_371_0_sva_dfm_1 = sigmoid_table_371_0_sva | (~ initialized_sva);
  assign sigmoid_table_372_0_sva_dfm_1 = sigmoid_table_372_0_sva | (~ initialized_sva);
  assign sigmoid_table_375_0_sva_dfm_1 = sigmoid_table_375_0_sva | (~ initialized_sva);
  assign sigmoid_table_376_0_sva_dfm_1 = sigmoid_table_376_0_sva | (~ initialized_sva);
  assign sigmoid_table_379_0_sva_dfm_1 = sigmoid_table_379_0_sva | (~ initialized_sva);
  assign sigmoid_table_380_0_sva_dfm_1 = sigmoid_table_380_0_sva | (~ initialized_sva);
  assign sigmoid_table_381_0_sva_dfm_1 = sigmoid_table_381_0_sva | (~ initialized_sva);
  assign sigmoid_table_385_0_sva_dfm_1 = sigmoid_table_385_0_sva | (~ initialized_sva);
  assign sigmoid_table_386_0_sva_dfm_1 = sigmoid_table_386_0_sva | (~ initialized_sva);
  assign sigmoid_table_387_0_sva_dfm_1 = sigmoid_table_387_0_sva | (~ initialized_sva);
  assign sigmoid_table_394_0_sva_dfm_1 = sigmoid_table_394_0_sva | (~ initialized_sva);
  assign sigmoid_table_395_0_sva_dfm_1 = sigmoid_table_395_0_sva | (~ initialized_sva);
  assign sigmoid_table_396_0_sva_dfm_1 = sigmoid_table_396_0_sva | (~ initialized_sva);
  assign sigmoid_table_397_0_sva_dfm_1 = sigmoid_table_397_0_sva | (~ initialized_sva);
  assign sigmoid_table_398_0_sva_dfm_1 = sigmoid_table_398_0_sva | (~ initialized_sva);
  assign sigmoid_table_399_0_sva_dfm_1 = sigmoid_table_399_0_sva | (~ initialized_sva);
  assign sigmoid_table_400_0_sva_dfm_1 = sigmoid_table_400_0_sva | (~ initialized_sva);
  assign sigmoid_table_401_0_sva_dfm_1 = sigmoid_table_401_0_sva | (~ initialized_sva);
  assign sigmoid_table_402_0_sva_dfm_1 = sigmoid_table_402_0_sva | (~ initialized_sva);
  assign sigmoid_table_403_0_sva_dfm_1 = sigmoid_table_403_0_sva | (~ initialized_sva);
  assign sigmoid_table_404_0_sva_dfm_1 = sigmoid_table_404_0_sva | (~ initialized_sva);
  assign sigmoid_table_405_0_sva_dfm_1 = sigmoid_table_405_0_sva | (~ initialized_sva);
  assign sigmoid_table_411_0_sva_dfm_1 = sigmoid_table_411_0_sva | (~ initialized_sva);
  assign sigmoid_table_412_0_sva_dfm_1 = sigmoid_table_412_0_sva | (~ initialized_sva);
  assign sigmoid_table_413_0_sva_dfm_1 = sigmoid_table_413_0_sva | (~ initialized_sva);
  assign sigmoid_table_417_0_sva_dfm_1 = sigmoid_table_417_0_sva | (~ initialized_sva);
  assign sigmoid_table_418_0_sva_dfm_1 = sigmoid_table_418_0_sva | (~ initialized_sva);
  assign sigmoid_table_421_0_sva_dfm_1 = sigmoid_table_421_0_sva | (~ initialized_sva);
  assign sigmoid_table_422_0_sva_dfm_1 = sigmoid_table_422_0_sva | (~ initialized_sva);
  assign sigmoid_table_425_0_sva_dfm_1 = sigmoid_table_425_0_sva | (~ initialized_sva);
  assign sigmoid_table_426_0_sva_dfm_1 = sigmoid_table_426_0_sva | (~ initialized_sva);
  assign sigmoid_table_428_0_sva_dfm_1 = sigmoid_table_428_0_sva | (~ initialized_sva);
  assign sigmoid_table_429_0_sva_dfm_1 = sigmoid_table_429_0_sva | (~ initialized_sva);
  assign sigmoid_table_431_0_sva_dfm_1 = sigmoid_table_431_0_sva | (~ initialized_sva);
  assign sigmoid_table_434_0_sva_dfm_1 = sigmoid_table_434_0_sva | (~ initialized_sva);
  assign sigmoid_table_436_0_sva_dfm_1 = sigmoid_table_436_0_sva | (~ initialized_sva);
  assign sigmoid_table_438_0_sva_dfm_1 = sigmoid_table_438_0_sva | (~ initialized_sva);
  assign sigmoid_table_441_0_sva_dfm_1 = sigmoid_table_441_0_sva | (~ initialized_sva);
  assign sigmoid_table_443_0_sva_dfm_1 = sigmoid_table_443_0_sva | (~ initialized_sva);
  assign sigmoid_table_446_0_sva_dfm_1 = sigmoid_table_446_0_sva | (~ initialized_sva);
  assign sigmoid_table_448_0_sva_dfm_1 = sigmoid_table_448_0_sva | (~ initialized_sva);
  assign sigmoid_table_450_0_sva_dfm_1 = sigmoid_table_450_0_sva | (~ initialized_sva);
  assign sigmoid_table_453_0_sva_dfm_1 = sigmoid_table_453_0_sva | (~ initialized_sva);
  assign sigmoid_table_455_0_sva_dfm_1 = sigmoid_table_455_0_sva | (~ initialized_sva);
  assign sigmoid_table_456_0_sva_dfm_1 = sigmoid_table_456_0_sva | (~ initialized_sva);
  assign sigmoid_table_458_0_sva_dfm_1 = sigmoid_table_458_0_sva | (~ initialized_sva);
  assign sigmoid_table_459_0_sva_dfm_1 = sigmoid_table_459_0_sva | (~ initialized_sva);
  assign sigmoid_table_462_0_sva_dfm_1 = sigmoid_table_462_0_sva | (~ initialized_sva);
  assign sigmoid_table_463_0_sva_dfm_1 = sigmoid_table_463_0_sva | (~ initialized_sva);
  assign sigmoid_table_466_0_sva_dfm_1 = sigmoid_table_466_0_sva | (~ initialized_sva);
  assign sigmoid_table_467_0_sva_dfm_1 = sigmoid_table_467_0_sva | (~ initialized_sva);
  assign sigmoid_table_470_0_sva_dfm_1 = sigmoid_table_470_0_sva | (~ initialized_sva);
  assign sigmoid_table_471_0_sva_dfm_1 = sigmoid_table_471_0_sva | (~ initialized_sva);
  assign sigmoid_table_472_0_sva_dfm_1 = sigmoid_table_472_0_sva | (~ initialized_sva);
  assign sigmoid_table_475_0_sva_dfm_1 = sigmoid_table_475_0_sva | (~ initialized_sva);
  assign sigmoid_table_476_0_sva_dfm_1 = sigmoid_table_476_0_sva | (~ initialized_sva);
  assign sigmoid_table_477_0_sva_dfm_1 = sigmoid_table_477_0_sva | (~ initialized_sva);
  assign sigmoid_table_478_0_sva_dfm_1 = sigmoid_table_478_0_sva | (~ initialized_sva);
  assign sigmoid_table_483_0_sva_dfm_1 = sigmoid_table_483_0_sva | (~ initialized_sva);
  assign sigmoid_table_484_0_sva_dfm_1 = sigmoid_table_484_0_sva | (~ initialized_sva);
  assign sigmoid_table_485_0_sva_dfm_1 = sigmoid_table_485_0_sva | (~ initialized_sva);
  assign sigmoid_table_486_0_sva_dfm_1 = sigmoid_table_486_0_sva | (~ initialized_sva);
  assign sigmoid_table_487_0_sva_dfm_1 = sigmoid_table_487_0_sva | (~ initialized_sva);
  assign sigmoid_table_488_0_sva_dfm_1 = sigmoid_table_488_0_sva | (~ initialized_sva);
  assign sigmoid_table_516_0_sva_dfm_1 = sigmoid_table_516_0_sva | (~ initialized_sva);
  assign sigmoid_table_517_0_sva_dfm_1 = sigmoid_table_517_0_sva | (~ initialized_sva);
  assign sigmoid_table_518_0_sva_dfm_1 = sigmoid_table_518_0_sva | (~ initialized_sva);
  assign sigmoid_table_519_0_sva_dfm_1 = sigmoid_table_519_0_sva | (~ initialized_sva);
  assign sigmoid_table_520_0_sva_dfm_1 = sigmoid_table_520_0_sva | (~ initialized_sva);
  assign sigmoid_table_521_0_sva_dfm_1 = sigmoid_table_521_0_sva | (~ initialized_sva);
  assign sigmoid_table_522_0_sva_dfm_1 = sigmoid_table_522_0_sva | (~ initialized_sva);
  assign sigmoid_table_523_0_sva_dfm_1 = sigmoid_table_523_0_sva | (~ initialized_sva);
  assign sigmoid_table_524_0_sva_dfm_1 = sigmoid_table_524_0_sva | (~ initialized_sva);
  assign sigmoid_table_525_0_sva_dfm_1 = sigmoid_table_525_0_sva | (~ initialized_sva);
  assign sigmoid_table_526_0_sva_dfm_1 = sigmoid_table_526_0_sva | (~ initialized_sva);
  assign sigmoid_table_527_0_sva_dfm_1 = sigmoid_table_527_0_sva | (~ initialized_sva);
  assign sigmoid_table_528_0_sva_dfm_1 = sigmoid_table_528_0_sva | (~ initialized_sva);
  assign sigmoid_table_529_0_sva_dfm_1 = sigmoid_table_529_0_sva | (~ initialized_sva);
  assign sigmoid_table_530_0_sva_dfm_1 = sigmoid_table_530_0_sva | (~ initialized_sva);
  assign sigmoid_table_531_0_sva_dfm_1 = sigmoid_table_531_0_sva | (~ initialized_sva);
  assign sigmoid_table_532_0_sva_dfm_1 = sigmoid_table_532_0_sva | (~ initialized_sva);
  assign sigmoid_table_533_0_sva_dfm_1 = sigmoid_table_533_0_sva | (~ initialized_sva);
  assign sigmoid_table_534_0_sva_dfm_1 = sigmoid_table_534_0_sva | (~ initialized_sva);
  assign sigmoid_table_535_0_sva_dfm_1 = sigmoid_table_535_0_sva | (~ initialized_sva);
  assign sigmoid_table_542_0_sva_dfm_1 = sigmoid_table_542_0_sva | (~ initialized_sva);
  assign sigmoid_table_543_0_sva_dfm_1 = sigmoid_table_543_0_sva | (~ initialized_sva);
  assign sigmoid_table_544_0_sva_dfm_1 = sigmoid_table_544_0_sva | (~ initialized_sva);
  assign sigmoid_table_545_0_sva_dfm_1 = sigmoid_table_545_0_sva | (~ initialized_sva);
  assign sigmoid_table_550_0_sva_dfm_1 = sigmoid_table_550_0_sva | (~ initialized_sva);
  assign sigmoid_table_551_0_sva_dfm_1 = sigmoid_table_551_0_sva | (~ initialized_sva);
  assign sigmoid_table_555_0_sva_dfm_1 = sigmoid_table_555_0_sva | (~ initialized_sva);
  assign sigmoid_table_556_0_sva_dfm_1 = sigmoid_table_556_0_sva | (~ initialized_sva);
  assign sigmoid_table_559_0_sva_dfm_1 = sigmoid_table_559_0_sva | (~ initialized_sva);
  assign sigmoid_table_560_0_sva_dfm_1 = sigmoid_table_560_0_sva | (~ initialized_sva);
  assign sigmoid_table_563_0_sva_dfm_1 = sigmoid_table_563_0_sva | (~ initialized_sva);
  assign sigmoid_table_564_0_sva_dfm_1 = sigmoid_table_564_0_sva | (~ initialized_sva);
  assign sigmoid_table_567_0_sva_dfm_1 = sigmoid_table_567_0_sva | (~ initialized_sva);
  assign sigmoid_table_570_0_sva_dfm_1 = sigmoid_table_570_0_sva | (~ initialized_sva);
  assign sigmoid_table_572_0_sva_dfm_1 = sigmoid_table_572_0_sva | (~ initialized_sva);
  assign sigmoid_table_573_0_sva_dfm_1 = sigmoid_table_573_0_sva | (~ initialized_sva);
  assign sigmoid_table_575_0_sva_dfm_1 = sigmoid_table_575_0_sva | (~ initialized_sva);
  assign sigmoid_table_577_0_sva_dfm_1 = sigmoid_table_577_0_sva | (~ initialized_sva);
  assign sigmoid_table_579_0_sva_dfm_1 = sigmoid_table_579_0_sva | (~ initialized_sva);
  assign sigmoid_table_580_0_sva_dfm_1 = sigmoid_table_580_0_sva | (~ initialized_sva);
  assign sigmoid_table_582_0_sva_dfm_1 = sigmoid_table_582_0_sva | (~ initialized_sva);
  assign sigmoid_table_584_0_sva_dfm_1 = sigmoid_table_584_0_sva | (~ initialized_sva);
  assign sigmoid_table_585_0_sva_dfm_1 = sigmoid_table_585_0_sva | (~ initialized_sva);
  assign sigmoid_table_587_0_sva_dfm_1 = sigmoid_table_587_0_sva | (~ initialized_sva);
  assign sigmoid_table_589_0_sva_dfm_1 = sigmoid_table_589_0_sva | (~ initialized_sva);
  assign sigmoid_table_591_0_sva_dfm_1 = sigmoid_table_591_0_sva | (~ initialized_sva);
  assign sigmoid_table_592_0_sva_dfm_1 = sigmoid_table_592_0_sva | (~ initialized_sva);
  assign sigmoid_table_594_0_sva_dfm_1 = sigmoid_table_594_0_sva | (~ initialized_sva);
  assign sigmoid_table_597_0_sva_dfm_1 = sigmoid_table_597_0_sva | (~ initialized_sva);
  assign sigmoid_table_600_0_sva_dfm_1 = sigmoid_table_600_0_sva | (~ initialized_sva);
  assign sigmoid_table_601_0_sva_dfm_1 = sigmoid_table_601_0_sva | (~ initialized_sva);
  assign sigmoid_table_604_0_sva_dfm_1 = sigmoid_table_604_0_sva | (~ initialized_sva);
  assign sigmoid_table_605_0_sva_dfm_1 = sigmoid_table_605_0_sva | (~ initialized_sva);
  assign sigmoid_table_608_0_sva_dfm_1 = sigmoid_table_608_0_sva | (~ initialized_sva);
  assign sigmoid_table_609_0_sva_dfm_1 = sigmoid_table_609_0_sva | (~ initialized_sva);
  assign sigmoid_table_610_0_sva_dfm_1 = sigmoid_table_610_0_sva | (~ initialized_sva);
  assign sigmoid_table_614_0_sva_dfm_1 = sigmoid_table_614_0_sva | (~ initialized_sva);
  assign sigmoid_table_615_0_sva_dfm_1 = sigmoid_table_615_0_sva | (~ initialized_sva);
  assign sigmoid_table_616_0_sva_dfm_1 = sigmoid_table_616_0_sva | (~ initialized_sva);
  assign sigmoid_table_617_0_sva_dfm_1 = sigmoid_table_617_0_sva | (~ initialized_sva);
  assign sigmoid_table_618_0_sva_dfm_1 = sigmoid_table_618_0_sva | (~ initialized_sva);
  assign sigmoid_table_631_0_sva_dfm_1 = sigmoid_table_631_0_sva | (~ initialized_sva);
  assign sigmoid_table_632_0_sva_dfm_1 = sigmoid_table_632_0_sva | (~ initialized_sva);
  assign sigmoid_table_633_0_sva_dfm_1 = sigmoid_table_633_0_sva | (~ initialized_sva);
  assign sigmoid_table_634_0_sva_dfm_1 = sigmoid_table_634_0_sva | (~ initialized_sva);
  assign sigmoid_table_635_0_sva_dfm_1 = sigmoid_table_635_0_sva | (~ initialized_sva);
  assign sigmoid_table_636_0_sva_dfm_1 = sigmoid_table_636_0_sva | (~ initialized_sva);
  assign sigmoid_table_640_0_sva_dfm_1 = sigmoid_table_640_0_sva | (~ initialized_sva);
  assign sigmoid_table_641_0_sva_dfm_1 = sigmoid_table_641_0_sva | (~ initialized_sva);
  assign sigmoid_table_642_0_sva_dfm_1 = sigmoid_table_642_0_sva | (~ initialized_sva);
  assign sigmoid_table_646_0_sva_dfm_1 = sigmoid_table_646_0_sva | (~ initialized_sva);
  assign sigmoid_table_647_0_sva_dfm_1 = sigmoid_table_647_0_sva | (~ initialized_sva);
  assign sigmoid_table_650_0_sva_dfm_1 = sigmoid_table_650_0_sva | (~ initialized_sva);
  assign sigmoid_table_651_0_sva_dfm_1 = sigmoid_table_651_0_sva | (~ initialized_sva);
  assign sigmoid_table_654_0_sva_dfm_1 = sigmoid_table_654_0_sva | (~ initialized_sva);
  assign sigmoid_table_657_0_sva_dfm_1 = sigmoid_table_657_0_sva | (~ initialized_sva);
  assign sigmoid_table_658_0_sva_dfm_1 = sigmoid_table_658_0_sva | (~ initialized_sva);
  assign sigmoid_table_660_0_sva_dfm_1 = sigmoid_table_660_0_sva | (~ initialized_sva);
  assign sigmoid_table_661_0_sva_dfm_1 = sigmoid_table_661_0_sva | (~ initialized_sva);
  assign sigmoid_table_663_0_sva_dfm_1 = sigmoid_table_663_0_sva | (~ initialized_sva);
  assign sigmoid_table_666_0_sva_dfm_1 = sigmoid_table_666_0_sva | (~ initialized_sva);
  assign sigmoid_table_668_0_sva_dfm_1 = sigmoid_table_668_0_sva | (~ initialized_sva);
  assign sigmoid_table_671_0_sva_dfm_1 = sigmoid_table_671_0_sva | (~ initialized_sva);
  assign sigmoid_table_673_0_sva_dfm_1 = sigmoid_table_673_0_sva | (~ initialized_sva);
  assign sigmoid_table_675_0_sva_dfm_1 = sigmoid_table_675_0_sva | (~ initialized_sva);
  assign sigmoid_table_677_0_sva_dfm_1 = sigmoid_table_677_0_sva | (~ initialized_sva);
  assign sigmoid_table_679_0_sva_dfm_1 = sigmoid_table_679_0_sva | (~ initialized_sva);
  assign sigmoid_table_681_0_sva_dfm_1 = sigmoid_table_681_0_sva | (~ initialized_sva);
  assign sigmoid_table_683_0_sva_dfm_1 = sigmoid_table_683_0_sva | (~ initialized_sva);
  assign sigmoid_table_685_0_sva_dfm_1 = sigmoid_table_685_0_sva | (~ initialized_sva);
  assign sigmoid_table_687_0_sva_dfm_1 = sigmoid_table_687_0_sva | (~ initialized_sva);
  assign sigmoid_table_689_0_sva_dfm_1 = sigmoid_table_689_0_sva | (~ initialized_sva);
  assign sigmoid_table_691_0_sva_dfm_1 = sigmoid_table_691_0_sva | (~ initialized_sva);
  assign sigmoid_table_692_0_sva_dfm_1 = sigmoid_table_692_0_sva | (~ initialized_sva);
  assign sigmoid_table_694_0_sva_dfm_1 = sigmoid_table_694_0_sva | (~ initialized_sva);
  assign sigmoid_table_696_0_sva_dfm_1 = sigmoid_table_696_0_sva | (~ initialized_sva);
  assign sigmoid_table_699_0_sva_dfm_1 = sigmoid_table_699_0_sva | (~ initialized_sva);
  assign sigmoid_table_701_0_sva_dfm_1 = sigmoid_table_701_0_sva | (~ initialized_sva);
  assign sigmoid_table_702_0_sva_dfm_1 = sigmoid_table_702_0_sva | (~ initialized_sva);
  assign sigmoid_table_704_0_sva_dfm_1 = sigmoid_table_704_0_sva | (~ initialized_sva);
  assign sigmoid_table_707_0_sva_dfm_1 = sigmoid_table_707_0_sva | (~ initialized_sva);
  assign sigmoid_table_710_0_sva_dfm_1 = sigmoid_table_710_0_sva | (~ initialized_sva);
  assign sigmoid_table_713_0_sva_dfm_1 = sigmoid_table_713_0_sva | (~ initialized_sva);
  assign sigmoid_table_716_0_sva_dfm_1 = sigmoid_table_716_0_sva | (~ initialized_sva);
  assign sigmoid_table_719_0_sva_dfm_1 = sigmoid_table_719_0_sva | (~ initialized_sva);
  assign sigmoid_table_720_0_sva_dfm_1 = sigmoid_table_720_0_sva | (~ initialized_sva);
  assign sigmoid_table_723_0_sva_dfm_1 = sigmoid_table_723_0_sva | (~ initialized_sva);
  assign sigmoid_table_726_0_sva_dfm_1 = sigmoid_table_726_0_sva | (~ initialized_sva);
  assign sigmoid_table_727_0_sva_dfm_1 = sigmoid_table_727_0_sva | (~ initialized_sva);
  assign sigmoid_table_730_0_sva_dfm_1 = sigmoid_table_730_0_sva | (~ initialized_sva);
  assign sigmoid_table_731_0_sva_dfm_1 = sigmoid_table_731_0_sva | (~ initialized_sva);
  assign sigmoid_table_734_0_sva_dfm_1 = sigmoid_table_734_0_sva | (~ initialized_sva);
  assign sigmoid_table_735_0_sva_dfm_1 = sigmoid_table_735_0_sva | (~ initialized_sva);
  assign sigmoid_table_736_0_sva_dfm_1 = sigmoid_table_736_0_sva | (~ initialized_sva);
  assign sigmoid_table_739_0_sva_dfm_1 = sigmoid_table_739_0_sva | (~ initialized_sva);
  assign sigmoid_table_740_0_sva_dfm_1 = sigmoid_table_740_0_sva | (~ initialized_sva);
  assign sigmoid_table_743_0_sva_dfm_1 = sigmoid_table_743_0_sva | (~ initialized_sva);
  assign sigmoid_table_744_0_sva_dfm_1 = sigmoid_table_744_0_sva | (~ initialized_sva);
  assign sigmoid_table_745_0_sva_dfm_1 = sigmoid_table_745_0_sva | (~ initialized_sva);
  assign sigmoid_table_748_0_sva_dfm_1 = sigmoid_table_748_0_sva | (~ initialized_sva);
  assign sigmoid_table_749_0_sva_dfm_1 = sigmoid_table_749_0_sva | (~ initialized_sva);
  assign sigmoid_table_750_0_sva_dfm_1 = sigmoid_table_750_0_sva | (~ initialized_sva);
  assign sigmoid_table_754_0_sva_dfm_1 = sigmoid_table_754_0_sva | (~ initialized_sva);
  assign sigmoid_table_755_0_sva_dfm_1 = sigmoid_table_755_0_sva | (~ initialized_sva);
  assign sigmoid_table_756_0_sva_dfm_1 = sigmoid_table_756_0_sva | (~ initialized_sva);
  assign sigmoid_table_760_0_sva_dfm_1 = sigmoid_table_760_0_sva | (~ initialized_sva);
  assign sigmoid_table_761_0_sva_dfm_1 = sigmoid_table_761_0_sva | (~ initialized_sva);
  assign sigmoid_table_762_0_sva_dfm_1 = sigmoid_table_762_0_sva | (~ initialized_sva);
  assign sigmoid_table_766_0_sva_dfm_1 = sigmoid_table_766_0_sva | (~ initialized_sva);
  assign sigmoid_table_767_0_sva_dfm_1 = sigmoid_table_767_0_sva | (~ initialized_sva);
  assign sigmoid_table_768_0_sva_dfm_1 = sigmoid_table_768_0_sva | (~ initialized_sva);
  assign sigmoid_table_769_0_sva_dfm_1 = sigmoid_table_769_0_sva | (~ initialized_sva);
  assign sigmoid_table_774_0_sva_dfm_1 = sigmoid_table_774_0_sva | (~ initialized_sva);
  assign sigmoid_table_775_0_sva_dfm_1 = sigmoid_table_775_0_sva | (~ initialized_sva);
  assign sigmoid_table_776_0_sva_dfm_1 = sigmoid_table_776_0_sva | (~ initialized_sva);
  assign sigmoid_table_777_0_sva_dfm_1 = sigmoid_table_777_0_sva | (~ initialized_sva);
  assign sigmoid_table_782_0_sva_dfm_1 = sigmoid_table_782_0_sva | (~ initialized_sva);
  assign sigmoid_table_783_0_sva_dfm_1 = sigmoid_table_783_0_sva | (~ initialized_sva);
  assign sigmoid_table_784_0_sva_dfm_1 = sigmoid_table_784_0_sva | (~ initialized_sva);
  assign sigmoid_table_785_0_sva_dfm_1 = sigmoid_table_785_0_sva | (~ initialized_sva);
  assign sigmoid_table_791_0_sva_dfm_1 = sigmoid_table_791_0_sva | (~ initialized_sva);
  assign sigmoid_table_792_0_sva_dfm_1 = sigmoid_table_792_0_sva | (~ initialized_sva);
  assign sigmoid_table_793_0_sva_dfm_1 = sigmoid_table_793_0_sva | (~ initialized_sva);
  assign sigmoid_table_794_0_sva_dfm_1 = sigmoid_table_794_0_sva | (~ initialized_sva);
  assign sigmoid_table_795_0_sva_dfm_1 = sigmoid_table_795_0_sva | (~ initialized_sva);
  assign sigmoid_table_802_0_sva_dfm_1 = sigmoid_table_802_0_sva | (~ initialized_sva);
  assign sigmoid_table_803_0_sva_dfm_1 = sigmoid_table_803_0_sva | (~ initialized_sva);
  assign sigmoid_table_804_0_sva_dfm_1 = sigmoid_table_804_0_sva | (~ initialized_sva);
  assign sigmoid_table_805_0_sva_dfm_1 = sigmoid_table_805_0_sva | (~ initialized_sva);
  assign sigmoid_table_806_0_sva_dfm_1 = sigmoid_table_806_0_sva | (~ initialized_sva);
  assign sigmoid_table_807_0_sva_dfm_1 = sigmoid_table_807_0_sva | (~ initialized_sva);
  assign sigmoid_table_815_0_sva_dfm_1 = sigmoid_table_815_0_sva | (~ initialized_sva);
  assign sigmoid_table_816_0_sva_dfm_1 = sigmoid_table_816_0_sva | (~ initialized_sva);
  assign sigmoid_table_817_0_sva_dfm_1 = sigmoid_table_817_0_sva | (~ initialized_sva);
  assign sigmoid_table_818_0_sva_dfm_1 = sigmoid_table_818_0_sva | (~ initialized_sva);
  assign sigmoid_table_819_0_sva_dfm_1 = sigmoid_table_819_0_sva | (~ initialized_sva);
  assign sigmoid_table_820_0_sva_dfm_1 = sigmoid_table_820_0_sva | (~ initialized_sva);
  assign sigmoid_table_821_0_sva_dfm_1 = sigmoid_table_821_0_sva | (~ initialized_sva);
  assign sigmoid_table_831_0_sva_dfm_1 = sigmoid_table_831_0_sva | (~ initialized_sva);
  assign sigmoid_table_832_0_sva_dfm_1 = sigmoid_table_832_0_sva | (~ initialized_sva);
  assign sigmoid_table_833_0_sva_dfm_1 = sigmoid_table_833_0_sva | (~ initialized_sva);
  assign sigmoid_table_834_0_sva_dfm_1 = sigmoid_table_834_0_sva | (~ initialized_sva);
  assign sigmoid_table_835_0_sva_dfm_1 = sigmoid_table_835_0_sva | (~ initialized_sva);
  assign sigmoid_table_836_0_sva_dfm_1 = sigmoid_table_836_0_sva | (~ initialized_sva);
  assign sigmoid_table_837_0_sva_dfm_1 = sigmoid_table_837_0_sva | (~ initialized_sva);
  assign sigmoid_table_838_0_sva_dfm_1 = sigmoid_table_838_0_sva | (~ initialized_sva);
  assign sigmoid_table_839_0_sva_dfm_1 = sigmoid_table_839_0_sva | (~ initialized_sva);
  assign sigmoid_table_840_0_sva_dfm_1 = sigmoid_table_840_0_sva | (~ initialized_sva);
  assign sigmoid_table_853_0_sva_dfm_1 = sigmoid_table_853_0_sva | (~ initialized_sva);
  assign sigmoid_table_854_0_sva_dfm_1 = sigmoid_table_854_0_sva | (~ initialized_sva);
  assign sigmoid_table_855_0_sva_dfm_1 = sigmoid_table_855_0_sva | (~ initialized_sva);
  assign sigmoid_table_856_0_sva_dfm_1 = sigmoid_table_856_0_sva | (~ initialized_sva);
  assign sigmoid_table_857_0_sva_dfm_1 = sigmoid_table_857_0_sva | (~ initialized_sva);
  assign sigmoid_table_858_0_sva_dfm_1 = sigmoid_table_858_0_sva | (~ initialized_sva);
  assign sigmoid_table_859_0_sva_dfm_1 = sigmoid_table_859_0_sva | (~ initialized_sva);
  assign sigmoid_table_860_0_sva_dfm_1 = sigmoid_table_860_0_sva | (~ initialized_sva);
  assign sigmoid_table_861_0_sva_dfm_1 = sigmoid_table_861_0_sva | (~ initialized_sva);
  assign sigmoid_table_862_0_sva_dfm_1 = sigmoid_table_862_0_sva | (~ initialized_sva);
  assign sigmoid_table_863_0_sva_dfm_1 = sigmoid_table_863_0_sva | (~ initialized_sva);
  assign sigmoid_table_864_0_sva_dfm_1 = sigmoid_table_864_0_sva | (~ initialized_sva);
  assign sigmoid_table_865_0_sva_dfm_1 = sigmoid_table_865_0_sva | (~ initialized_sva);
  assign sigmoid_table_866_0_sva_dfm_1 = sigmoid_table_866_0_sva | (~ initialized_sva);
  assign sigmoid_table_885_0_sva_dfm_1 = sigmoid_table_885_0_sva | (~ initialized_sva);
  assign sigmoid_table_886_0_sva_dfm_1 = sigmoid_table_886_0_sva | (~ initialized_sva);
  assign sigmoid_table_887_0_sva_dfm_1 = sigmoid_table_887_0_sva | (~ initialized_sva);
  assign sigmoid_table_888_0_sva_dfm_1 = sigmoid_table_888_0_sva | (~ initialized_sva);
  assign sigmoid_table_889_0_sva_dfm_1 = sigmoid_table_889_0_sva | (~ initialized_sva);
  assign sigmoid_table_890_0_sva_dfm_1 = sigmoid_table_890_0_sva | (~ initialized_sva);
  assign sigmoid_table_891_0_sva_dfm_1 = sigmoid_table_891_0_sva | (~ initialized_sva);
  assign sigmoid_table_892_0_sva_dfm_1 = sigmoid_table_892_0_sva | (~ initialized_sva);
  assign sigmoid_table_893_0_sva_dfm_1 = sigmoid_table_893_0_sva | (~ initialized_sva);
  assign sigmoid_table_894_0_sva_dfm_1 = sigmoid_table_894_0_sva | (~ initialized_sva);
  assign sigmoid_table_895_0_sva_dfm_1 = sigmoid_table_895_0_sva | (~ initialized_sva);
  assign sigmoid_table_896_0_sva_dfm_1 = sigmoid_table_896_0_sva | (~ initialized_sva);
  assign sigmoid_table_897_0_sva_dfm_1 = sigmoid_table_897_0_sva | (~ initialized_sva);
  assign sigmoid_table_898_0_sva_dfm_1 = sigmoid_table_898_0_sva | (~ initialized_sva);
  assign sigmoid_table_899_0_sva_dfm_1 = sigmoid_table_899_0_sva | (~ initialized_sva);
  assign sigmoid_table_900_0_sva_dfm_1 = sigmoid_table_900_0_sva | (~ initialized_sva);
  assign sigmoid_table_901_0_sva_dfm_1 = sigmoid_table_901_0_sva | (~ initialized_sva);
  assign sigmoid_table_902_0_sva_dfm_1 = sigmoid_table_902_0_sva | (~ initialized_sva);
  assign sigmoid_table_903_0_sva_dfm_1 = sigmoid_table_903_0_sva | (~ initialized_sva);
  assign sigmoid_table_904_0_sva_dfm_1 = sigmoid_table_904_0_sva | (~ initialized_sva);
  assign sigmoid_table_905_0_sva_dfm_1 = sigmoid_table_905_0_sva | (~ initialized_sva);
  assign sigmoid_table_906_0_sva_dfm_1 = sigmoid_table_906_0_sva | (~ initialized_sva);
  assign sigmoid_table_907_0_sva_dfm_1 = sigmoid_table_907_0_sva | (~ initialized_sva);
  assign sigmoid_table_908_0_sva_dfm_1 = sigmoid_table_908_0_sva | (~ initialized_sva);
  assign sigmoid_table_909_0_sva_dfm_1 = sigmoid_table_909_0_sva | (~ initialized_sva);
  assign sigmoid_table_910_0_sva_dfm_1 = sigmoid_table_910_0_sva | (~ initialized_sva);
  assign sigmoid_table_955_0_sva_dfm_1 = sigmoid_table_955_0_sva | (~ initialized_sva);
  assign sigmoid_table_956_0_sva_dfm_1 = sigmoid_table_956_0_sva | (~ initialized_sva);
  assign sigmoid_table_957_0_sva_dfm_1 = sigmoid_table_957_0_sva | (~ initialized_sva);
  assign sigmoid_table_958_0_sva_dfm_1 = sigmoid_table_958_0_sva | (~ initialized_sva);
  assign sigmoid_table_959_0_sva_dfm_1 = sigmoid_table_959_0_sva | (~ initialized_sva);
  assign sigmoid_table_960_0_sva_dfm_1 = sigmoid_table_960_0_sva | (~ initialized_sva);
  assign sigmoid_table_961_0_sva_dfm_1 = sigmoid_table_961_0_sva | (~ initialized_sva);
  assign sigmoid_table_962_0_sva_dfm_1 = sigmoid_table_962_0_sva | (~ initialized_sva);
  assign sigmoid_table_963_0_sva_dfm_1 = sigmoid_table_963_0_sva | (~ initialized_sva);
  assign sigmoid_table_964_0_sva_dfm_1 = sigmoid_table_964_0_sva | (~ initialized_sva);
  assign sigmoid_table_965_0_sva_dfm_1 = sigmoid_table_965_0_sva | (~ initialized_sva);
  assign sigmoid_table_966_0_sva_dfm_1 = sigmoid_table_966_0_sva | (~ initialized_sva);
  assign sigmoid_table_967_0_sva_dfm_1 = sigmoid_table_967_0_sva | (~ initialized_sva);
  assign sigmoid_table_968_0_sva_dfm_1 = sigmoid_table_968_0_sva | (~ initialized_sva);
  assign sigmoid_table_969_0_sva_dfm_1 = sigmoid_table_969_0_sva | (~ initialized_sva);
  assign sigmoid_table_970_0_sva_dfm_1 = sigmoid_table_970_0_sva | (~ initialized_sva);
  assign sigmoid_table_971_0_sva_dfm_1 = sigmoid_table_971_0_sva | (~ initialized_sva);
  assign sigmoid_table_972_0_sva_dfm_1 = sigmoid_table_972_0_sva | (~ initialized_sva);
  assign sigmoid_table_973_0_sva_dfm_1 = sigmoid_table_973_0_sva | (~ initialized_sva);
  assign sigmoid_table_974_0_sva_dfm_1 = sigmoid_table_974_0_sva | (~ initialized_sva);
  assign sigmoid_table_975_0_sva_dfm_1 = sigmoid_table_975_0_sva | (~ initialized_sva);
  assign sigmoid_table_976_0_sva_dfm_1 = sigmoid_table_976_0_sva | (~ initialized_sva);
  assign sigmoid_table_977_0_sva_dfm_1 = sigmoid_table_977_0_sva | (~ initialized_sva);
  assign sigmoid_table_978_0_sva_dfm_1 = sigmoid_table_978_0_sva | (~ initialized_sva);
  assign sigmoid_table_979_0_sva_dfm_1 = sigmoid_table_979_0_sva | (~ initialized_sva);
  assign sigmoid_table_980_0_sva_dfm_1 = sigmoid_table_980_0_sva | (~ initialized_sva);
  assign sigmoid_table_981_0_sva_dfm_1 = sigmoid_table_981_0_sva | (~ initialized_sva);
  assign sigmoid_table_982_0_sva_dfm_1 = sigmoid_table_982_0_sva | (~ initialized_sva);
  assign sigmoid_table_983_0_sva_dfm_1 = sigmoid_table_983_0_sva | (~ initialized_sva);
  assign sigmoid_table_984_0_sva_dfm_1 = sigmoid_table_984_0_sva | (~ initialized_sva);
  assign sigmoid_table_985_0_sva_dfm_1 = sigmoid_table_985_0_sva | (~ initialized_sva);
  assign sigmoid_table_986_0_sva_dfm_1 = sigmoid_table_986_0_sva | (~ initialized_sva);
  assign sigmoid_table_987_0_sva_dfm_1 = sigmoid_table_987_0_sva | (~ initialized_sva);
  assign sigmoid_table_988_0_sva_dfm_1 = sigmoid_table_988_0_sva | (~ initialized_sva);
  assign sigmoid_table_989_0_sva_dfm_1 = sigmoid_table_989_0_sva | (~ initialized_sva);
  assign sigmoid_table_990_0_sva_dfm_1 = sigmoid_table_990_0_sva | (~ initialized_sva);
  assign sigmoid_table_991_0_sva_dfm_1 = sigmoid_table_991_0_sva | (~ initialized_sva);
  assign sigmoid_table_992_0_sva_dfm_1 = sigmoid_table_992_0_sva | (~ initialized_sva);
  assign sigmoid_table_993_0_sva_dfm_1 = sigmoid_table_993_0_sva | (~ initialized_sva);
  assign sigmoid_table_994_0_sva_dfm_1 = sigmoid_table_994_0_sva | (~ initialized_sva);
  assign sigmoid_table_995_0_sva_dfm_1 = sigmoid_table_995_0_sva | (~ initialized_sva);
  assign sigmoid_table_996_0_sva_dfm_1 = sigmoid_table_996_0_sva | (~ initialized_sva);
  assign sigmoid_table_997_0_sva_dfm_1 = sigmoid_table_997_0_sva | (~ initialized_sva);
  assign sigmoid_table_998_0_sva_dfm_1 = sigmoid_table_998_0_sva | (~ initialized_sva);
  assign sigmoid_table_999_0_sva_dfm_1 = sigmoid_table_999_0_sva | (~ initialized_sva);
  assign sigmoid_table_1000_0_sva_dfm_1 = sigmoid_table_1000_0_sva | (~ initialized_sva);
  assign sigmoid_table_1001_0_sva_dfm_1 = sigmoid_table_1001_0_sva | (~ initialized_sva);
  assign sigmoid_table_1002_0_sva_dfm_1 = sigmoid_table_1002_0_sva | (~ initialized_sva);
  assign sigmoid_table_1003_0_sva_dfm_1 = sigmoid_table_1003_0_sva | (~ initialized_sva);
  assign sigmoid_table_1004_0_sva_dfm_1 = sigmoid_table_1004_0_sva | (~ initialized_sva);
  assign sigmoid_table_1005_0_sva_dfm_1 = sigmoid_table_1005_0_sva | (~ initialized_sva);
  assign sigmoid_table_1006_0_sva_dfm_1 = sigmoid_table_1006_0_sva | (~ initialized_sva);
  assign sigmoid_table_1007_0_sva_dfm_1 = sigmoid_table_1007_0_sva | (~ initialized_sva);
  assign sigmoid_table_1008_0_sva_dfm_1 = sigmoid_table_1008_0_sva | (~ initialized_sva);
  assign sigmoid_table_1009_0_sva_dfm_1 = sigmoid_table_1009_0_sva | (~ initialized_sva);
  assign sigmoid_table_1010_0_sva_dfm_1 = sigmoid_table_1010_0_sva | (~ initialized_sva);
  assign sigmoid_table_1011_0_sva_dfm_1 = sigmoid_table_1011_0_sva | (~ initialized_sva);
  assign sigmoid_table_1012_0_sva_dfm_1 = sigmoid_table_1012_0_sva | (~ initialized_sva);
  assign sigmoid_table_1013_0_sva_dfm_1 = sigmoid_table_1013_0_sva | (~ initialized_sva);
  assign sigmoid_table_1014_0_sva_dfm_1 = sigmoid_table_1014_0_sva | (~ initialized_sva);
  assign sigmoid_table_1015_0_sva_dfm_1 = sigmoid_table_1015_0_sva | (~ initialized_sva);
  assign sigmoid_table_1016_0_sva_dfm_1 = sigmoid_table_1016_0_sva | (~ initialized_sva);
  assign sigmoid_table_1017_0_sva_dfm_1 = sigmoid_table_1017_0_sva | (~ initialized_sva);
  assign sigmoid_table_1018_0_sva_dfm_1 = sigmoid_table_1018_0_sva | (~ initialized_sva);
  assign sigmoid_table_1019_0_sva_dfm_1 = sigmoid_table_1019_0_sva | (~ initialized_sva);
  assign sigmoid_table_1020_0_sva_dfm_1 = sigmoid_table_1020_0_sva | (~ initialized_sva);
  assign sigmoid_table_1021_0_sva_dfm_1 = sigmoid_table_1021_0_sva | (~ initialized_sva);
  assign sigmoid_table_1022_0_sva_dfm_1 = sigmoid_table_1022_0_sva | (~ initialized_sva);
  assign sigmoid_table_1023_0_sva_dfm_1 = sigmoid_table_1023_0_sva | (~ initialized_sva);
  assign sigmoid_table_512_9_sva_dfm_1 = sigmoid_table_512_9_sva | (~ initialized_sva);
  assign sigmoid_table_513_9_sva_dfm_1 = sigmoid_table_513_9_sva | (~ initialized_sva);
  assign sigmoid_table_514_9_sva_dfm_1 = sigmoid_table_514_9_sva | (~ initialized_sva);
  assign sigmoid_table_515_9_sva_dfm_1 = sigmoid_table_515_9_sva | (~ initialized_sva);
  assign sigmoid_table_516_9_sva_dfm_1 = sigmoid_table_516_9_sva | (~ initialized_sva);
  assign sigmoid_table_517_9_sva_dfm_1 = sigmoid_table_517_9_sva | (~ initialized_sva);
  assign sigmoid_table_518_9_sva_dfm_1 = sigmoid_table_518_9_sva | (~ initialized_sva);
  assign sigmoid_table_519_9_sva_dfm_1 = sigmoid_table_519_9_sva | (~ initialized_sva);
  assign sigmoid_table_520_9_sva_dfm_1 = sigmoid_table_520_9_sva | (~ initialized_sva);
  assign sigmoid_table_521_9_sva_dfm_1 = sigmoid_table_521_9_sva | (~ initialized_sva);
  assign sigmoid_table_522_9_sva_dfm_1 = sigmoid_table_522_9_sva | (~ initialized_sva);
  assign sigmoid_table_523_9_sva_dfm_1 = sigmoid_table_523_9_sva | (~ initialized_sva);
  assign sigmoid_table_524_9_sva_dfm_1 = sigmoid_table_524_9_sva | (~ initialized_sva);
  assign sigmoid_table_525_9_sva_dfm_1 = sigmoid_table_525_9_sva | (~ initialized_sva);
  assign sigmoid_table_526_9_sva_dfm_1 = sigmoid_table_526_9_sva | (~ initialized_sva);
  assign sigmoid_table_527_9_sva_dfm_1 = sigmoid_table_527_9_sva | (~ initialized_sva);
  assign sigmoid_table_528_9_sva_dfm_1 = sigmoid_table_528_9_sva | (~ initialized_sva);
  assign sigmoid_table_529_9_sva_dfm_1 = sigmoid_table_529_9_sva | (~ initialized_sva);
  assign sigmoid_table_530_9_sva_dfm_1 = sigmoid_table_530_9_sva | (~ initialized_sva);
  assign sigmoid_table_531_9_sva_dfm_1 = sigmoid_table_531_9_sva | (~ initialized_sva);
  assign sigmoid_table_532_9_sva_dfm_1 = sigmoid_table_532_9_sva | (~ initialized_sva);
  assign sigmoid_table_533_9_sva_dfm_1 = sigmoid_table_533_9_sva | (~ initialized_sva);
  assign sigmoid_table_534_9_sva_dfm_1 = sigmoid_table_534_9_sva | (~ initialized_sva);
  assign sigmoid_table_535_9_sva_dfm_1 = sigmoid_table_535_9_sva | (~ initialized_sva);
  assign sigmoid_table_536_9_sva_dfm_1 = sigmoid_table_536_9_sva | (~ initialized_sva);
  assign sigmoid_table_537_9_sva_dfm_1 = sigmoid_table_537_9_sva | (~ initialized_sva);
  assign sigmoid_table_538_9_sva_dfm_1 = sigmoid_table_538_9_sva | (~ initialized_sva);
  assign sigmoid_table_539_9_sva_dfm_1 = sigmoid_table_539_9_sva | (~ initialized_sva);
  assign sigmoid_table_540_9_sva_dfm_1 = sigmoid_table_540_9_sva | (~ initialized_sva);
  assign sigmoid_table_541_9_sva_dfm_1 = sigmoid_table_541_9_sva | (~ initialized_sva);
  assign sigmoid_table_542_9_sva_dfm_1 = sigmoid_table_542_9_sva | (~ initialized_sva);
  assign sigmoid_table_543_9_sva_dfm_1 = sigmoid_table_543_9_sva | (~ initialized_sva);
  assign sigmoid_table_544_9_sva_dfm_1 = sigmoid_table_544_9_sva | (~ initialized_sva);
  assign sigmoid_table_545_9_sva_dfm_1 = sigmoid_table_545_9_sva | (~ initialized_sva);
  assign sigmoid_table_546_9_sva_dfm_1 = sigmoid_table_546_9_sva | (~ initialized_sva);
  assign sigmoid_table_547_9_sva_dfm_1 = sigmoid_table_547_9_sva | (~ initialized_sva);
  assign sigmoid_table_548_9_sva_dfm_1 = sigmoid_table_548_9_sva | (~ initialized_sva);
  assign sigmoid_table_549_9_sva_dfm_1 = sigmoid_table_549_9_sva | (~ initialized_sva);
  assign sigmoid_table_550_9_sva_dfm_1 = sigmoid_table_550_9_sva | (~ initialized_sva);
  assign sigmoid_table_551_9_sva_dfm_1 = sigmoid_table_551_9_sva | (~ initialized_sva);
  assign sigmoid_table_552_9_sva_dfm_1 = sigmoid_table_552_9_sva | (~ initialized_sva);
  assign sigmoid_table_553_9_sva_dfm_1 = sigmoid_table_553_9_sva | (~ initialized_sva);
  assign sigmoid_table_554_9_sva_dfm_1 = sigmoid_table_554_9_sva | (~ initialized_sva);
  assign sigmoid_table_555_9_sva_dfm_1 = sigmoid_table_555_9_sva | (~ initialized_sva);
  assign sigmoid_table_556_9_sva_dfm_1 = sigmoid_table_556_9_sva | (~ initialized_sva);
  assign sigmoid_table_557_9_sva_dfm_1 = sigmoid_table_557_9_sva | (~ initialized_sva);
  assign sigmoid_table_558_9_sva_dfm_1 = sigmoid_table_558_9_sva | (~ initialized_sva);
  assign sigmoid_table_559_9_sva_dfm_1 = sigmoid_table_559_9_sva | (~ initialized_sva);
  assign sigmoid_table_560_9_sva_dfm_1 = sigmoid_table_560_9_sva | (~ initialized_sva);
  assign sigmoid_table_561_9_sva_dfm_1 = sigmoid_table_561_9_sva | (~ initialized_sva);
  assign sigmoid_table_562_9_sva_dfm_1 = sigmoid_table_562_9_sva | (~ initialized_sva);
  assign sigmoid_table_563_9_sva_dfm_1 = sigmoid_table_563_9_sva | (~ initialized_sva);
  assign sigmoid_table_564_9_sva_dfm_1 = sigmoid_table_564_9_sva | (~ initialized_sva);
  assign sigmoid_table_565_9_sva_dfm_1 = sigmoid_table_565_9_sva | (~ initialized_sva);
  assign sigmoid_table_566_9_sva_dfm_1 = sigmoid_table_566_9_sva | (~ initialized_sva);
  assign sigmoid_table_567_9_sva_dfm_1 = sigmoid_table_567_9_sva | (~ initialized_sva);
  assign sigmoid_table_568_9_sva_dfm_1 = sigmoid_table_568_9_sva | (~ initialized_sva);
  assign sigmoid_table_569_9_sva_dfm_1 = sigmoid_table_569_9_sva | (~ initialized_sva);
  assign sigmoid_table_570_9_sva_dfm_1 = sigmoid_table_570_9_sva | (~ initialized_sva);
  assign sigmoid_table_571_9_sva_dfm_1 = sigmoid_table_571_9_sva | (~ initialized_sva);
  assign sigmoid_table_572_9_sva_dfm_1 = sigmoid_table_572_9_sva | (~ initialized_sva);
  assign sigmoid_table_573_9_sva_dfm_1 = sigmoid_table_573_9_sva | (~ initialized_sva);
  assign sigmoid_table_574_9_sva_dfm_1 = sigmoid_table_574_9_sva | (~ initialized_sva);
  assign sigmoid_table_575_9_sva_dfm_1 = sigmoid_table_575_9_sva | (~ initialized_sva);
  assign sigmoid_table_576_9_sva_dfm_1 = sigmoid_table_576_9_sva | (~ initialized_sva);
  assign sigmoid_table_577_9_sva_dfm_1 = sigmoid_table_577_9_sva | (~ initialized_sva);
  assign sigmoid_table_578_9_sva_dfm_1 = sigmoid_table_578_9_sva | (~ initialized_sva);
  assign sigmoid_table_579_9_sva_dfm_1 = sigmoid_table_579_9_sva | (~ initialized_sva);
  assign sigmoid_table_580_9_sva_dfm_1 = sigmoid_table_580_9_sva | (~ initialized_sva);
  assign sigmoid_table_581_9_sva_dfm_1 = sigmoid_table_581_9_sva | (~ initialized_sva);
  assign sigmoid_table_582_9_sva_dfm_1 = sigmoid_table_582_9_sva | (~ initialized_sva);
  assign sigmoid_table_583_8_sva_dfm_1 = sigmoid_table_583_8_sva | (~ initialized_sva);
  assign sigmoid_table_584_8_sva_dfm_1 = sigmoid_table_584_8_sva | (~ initialized_sva);
  assign sigmoid_table_585_8_sva_dfm_1 = sigmoid_table_585_8_sva | (~ initialized_sva);
  assign sigmoid_table_586_8_sva_dfm_1 = sigmoid_table_586_8_sva | (~ initialized_sva);
  assign sigmoid_table_587_8_sva_dfm_1 = sigmoid_table_587_8_sva | (~ initialized_sva);
  assign sigmoid_table_588_8_sva_dfm_1 = sigmoid_table_588_8_sva | (~ initialized_sva);
  assign sigmoid_table_589_8_sva_dfm_1 = sigmoid_table_589_8_sva | (~ initialized_sva);
  assign sigmoid_table_590_8_sva_dfm_1 = sigmoid_table_590_8_sva | (~ initialized_sva);
  assign sigmoid_table_591_8_sva_dfm_1 = sigmoid_table_591_8_sva | (~ initialized_sva);
  assign sigmoid_table_592_8_sva_dfm_1 = sigmoid_table_592_8_sva | (~ initialized_sva);
  assign sigmoid_table_593_8_sva_dfm_1 = sigmoid_table_593_8_sva | (~ initialized_sva);
  assign sigmoid_table_594_8_sva_dfm_1 = sigmoid_table_594_8_sva | (~ initialized_sva);
  assign sigmoid_table_595_8_sva_dfm_1 = sigmoid_table_595_8_sva | (~ initialized_sva);
  assign sigmoid_table_596_8_sva_dfm_1 = sigmoid_table_596_8_sva | (~ initialized_sva);
  assign sigmoid_table_597_8_sva_dfm_1 = sigmoid_table_597_8_sva | (~ initialized_sva);
  assign sigmoid_table_598_8_sva_dfm_1 = sigmoid_table_598_8_sva | (~ initialized_sva);
  assign sigmoid_table_599_8_sva_dfm_1 = sigmoid_table_599_8_sva | (~ initialized_sva);
  assign sigmoid_table_600_8_sva_dfm_1 = sigmoid_table_600_8_sva | (~ initialized_sva);
  assign sigmoid_table_601_8_sva_dfm_1 = sigmoid_table_601_8_sva | (~ initialized_sva);
  assign sigmoid_table_602_8_sva_dfm_1 = sigmoid_table_602_8_sva | (~ initialized_sva);
  assign sigmoid_table_603_8_sva_dfm_1 = sigmoid_table_603_8_sva | (~ initialized_sva);
  assign sigmoid_table_604_8_sva_dfm_1 = sigmoid_table_604_8_sva | (~ initialized_sva);
  assign sigmoid_table_605_8_sva_dfm_1 = sigmoid_table_605_8_sva | (~ initialized_sva);
  assign sigmoid_table_606_8_sva_dfm_1 = sigmoid_table_606_8_sva | (~ initialized_sva);
  assign sigmoid_table_607_8_sva_dfm_1 = sigmoid_table_607_8_sva | (~ initialized_sva);
  assign sigmoid_table_608_8_sva_dfm_1 = sigmoid_table_608_8_sva | (~ initialized_sva);
  assign sigmoid_table_609_8_sva_dfm_1 = sigmoid_table_609_8_sva | (~ initialized_sva);
  assign sigmoid_table_610_8_sva_dfm_1 = sigmoid_table_610_8_sva | (~ initialized_sva);
  assign sigmoid_table_611_8_sva_dfm_1 = sigmoid_table_611_8_sva | (~ initialized_sva);
  assign sigmoid_table_612_8_sva_dfm_1 = sigmoid_table_612_8_sva | (~ initialized_sva);
  assign sigmoid_table_613_8_sva_dfm_1 = sigmoid_table_613_8_sva | (~ initialized_sva);
  assign sigmoid_table_614_8_sva_dfm_1 = sigmoid_table_614_8_sva | (~ initialized_sva);
  assign sigmoid_table_615_8_sva_dfm_1 = sigmoid_table_615_8_sva | (~ initialized_sva);
  assign sigmoid_table_616_8_sva_dfm_1 = sigmoid_table_616_8_sva | (~ initialized_sva);
  assign sigmoid_table_617_8_sva_dfm_1 = sigmoid_table_617_8_sva | (~ initialized_sva);
  assign sigmoid_table_618_8_sva_dfm_1 = sigmoid_table_618_8_sva | (~ initialized_sva);
  assign sigmoid_table_619_8_sva_dfm_1 = sigmoid_table_619_8_sva | (~ initialized_sva);
  assign sigmoid_table_620_8_sva_dfm_1 = sigmoid_table_620_8_sva | (~ initialized_sva);
  assign sigmoid_table_621_8_sva_dfm_1 = sigmoid_table_621_8_sva | (~ initialized_sva);
  assign sigmoid_table_622_8_sva_dfm_1 = sigmoid_table_622_8_sva | (~ initialized_sva);
  assign sigmoid_table_623_8_sva_dfm_1 = sigmoid_table_623_8_sva | (~ initialized_sva);
  assign sigmoid_table_624_8_sva_dfm_1 = sigmoid_table_624_8_sva | (~ initialized_sva);
  assign sigmoid_table_625_8_sva_dfm_1 = sigmoid_table_625_8_sva | (~ initialized_sva);
  assign sigmoid_table_626_8_sva_dfm_1 = sigmoid_table_626_8_sva | (~ initialized_sva);
  assign sigmoid_table_627_8_sva_dfm_1 = sigmoid_table_627_8_sva | (~ initialized_sva);
  assign sigmoid_table_628_8_sva_dfm_1 = sigmoid_table_628_8_sva | (~ initialized_sva);
  assign sigmoid_table_629_8_sva_dfm_1 = sigmoid_table_629_8_sva | (~ initialized_sva);
  assign sigmoid_table_630_8_sva_dfm_1 = sigmoid_table_630_8_sva | (~ initialized_sva);
  assign sigmoid_table_631_8_sva_dfm_1 = sigmoid_table_631_8_sva | (~ initialized_sva);
  assign sigmoid_table_632_8_sva_dfm_1 = sigmoid_table_632_8_sva | (~ initialized_sva);
  assign sigmoid_table_633_8_sva_dfm_1 = sigmoid_table_633_8_sva | (~ initialized_sva);
  assign sigmoid_table_634_8_sva_dfm_1 = sigmoid_table_634_8_sva | (~ initialized_sva);
  assign sigmoid_table_635_8_sva_dfm_1 = sigmoid_table_635_8_sva | (~ initialized_sva);
  assign sigmoid_table_636_8_sva_dfm_1 = sigmoid_table_636_8_sva | (~ initialized_sva);
  assign sigmoid_table_637_7_sva_dfm_1 = sigmoid_table_637_7_sva | (~ initialized_sva);
  assign sigmoid_table_638_7_sva_dfm_1 = sigmoid_table_638_7_sva | (~ initialized_sva);
  assign sigmoid_table_639_7_sva_dfm_1 = sigmoid_table_639_7_sva | (~ initialized_sva);
  assign sigmoid_table_640_7_sva_dfm_1 = sigmoid_table_640_7_sva | (~ initialized_sva);
  assign sigmoid_table_641_7_sva_dfm_1 = sigmoid_table_641_7_sva | (~ initialized_sva);
  assign sigmoid_table_642_7_sva_dfm_1 = sigmoid_table_642_7_sva | (~ initialized_sva);
  assign sigmoid_table_643_7_sva_dfm_1 = sigmoid_table_643_7_sva | (~ initialized_sva);
  assign sigmoid_table_644_7_sva_dfm_1 = sigmoid_table_644_7_sva | (~ initialized_sva);
  assign sigmoid_table_645_7_sva_dfm_1 = sigmoid_table_645_7_sva | (~ initialized_sva);
  assign sigmoid_table_646_7_sva_dfm_1 = sigmoid_table_646_7_sva | (~ initialized_sva);
  assign sigmoid_table_647_7_sva_dfm_1 = sigmoid_table_647_7_sva | (~ initialized_sva);
  assign sigmoid_table_648_7_sva_dfm_1 = sigmoid_table_648_7_sva | (~ initialized_sva);
  assign sigmoid_table_649_7_sva_dfm_1 = sigmoid_table_649_7_sva | (~ initialized_sva);
  assign sigmoid_table_650_7_sva_dfm_1 = sigmoid_table_650_7_sva | (~ initialized_sva);
  assign sigmoid_table_651_7_sva_dfm_1 = sigmoid_table_651_7_sva | (~ initialized_sva);
  assign sigmoid_table_652_7_sva_dfm_1 = sigmoid_table_652_7_sva | (~ initialized_sva);
  assign sigmoid_table_653_7_sva_dfm_1 = sigmoid_table_653_7_sva | (~ initialized_sva);
  assign sigmoid_table_654_7_sva_dfm_1 = sigmoid_table_654_7_sva | (~ initialized_sva);
  assign sigmoid_table_655_7_sva_dfm_1 = sigmoid_table_655_7_sva | (~ initialized_sva);
  assign sigmoid_table_656_7_sva_dfm_1 = sigmoid_table_656_7_sva | (~ initialized_sva);
  assign sigmoid_table_657_7_sva_dfm_1 = sigmoid_table_657_7_sva | (~ initialized_sva);
  assign sigmoid_table_658_7_sva_dfm_1 = sigmoid_table_658_7_sva | (~ initialized_sva);
  assign sigmoid_table_659_7_sva_dfm_1 = sigmoid_table_659_7_sva | (~ initialized_sva);
  assign sigmoid_table_660_7_sva_dfm_1 = sigmoid_table_660_7_sva | (~ initialized_sva);
  assign sigmoid_table_661_7_sva_dfm_1 = sigmoid_table_661_7_sva | (~ initialized_sva);
  assign sigmoid_table_662_7_sva_dfm_1 = sigmoid_table_662_7_sva | (~ initialized_sva);
  assign sigmoid_table_663_7_sva_dfm_1 = sigmoid_table_663_7_sva | (~ initialized_sva);
  assign sigmoid_table_664_7_sva_dfm_1 = sigmoid_table_664_7_sva | (~ initialized_sva);
  assign sigmoid_table_665_7_sva_dfm_1 = sigmoid_table_665_7_sva | (~ initialized_sva);
  assign sigmoid_table_666_7_sva_dfm_1 = sigmoid_table_666_7_sva | (~ initialized_sva);
  assign sigmoid_table_667_7_sva_dfm_1 = sigmoid_table_667_7_sva | (~ initialized_sva);
  assign sigmoid_table_668_7_sva_dfm_1 = sigmoid_table_668_7_sva | (~ initialized_sva);
  assign sigmoid_table_669_7_sva_dfm_1 = sigmoid_table_669_7_sva | (~ initialized_sva);
  assign sigmoid_table_670_7_sva_dfm_1 = sigmoid_table_670_7_sva | (~ initialized_sva);
  assign sigmoid_table_671_7_sva_dfm_1 = sigmoid_table_671_7_sva | (~ initialized_sva);
  assign sigmoid_table_672_7_sva_dfm_1 = sigmoid_table_672_7_sva | (~ initialized_sva);
  assign sigmoid_table_673_7_sva_dfm_1 = sigmoid_table_673_7_sva | (~ initialized_sva);
  assign sigmoid_table_674_7_sva_dfm_1 = sigmoid_table_674_7_sva | (~ initialized_sva);
  assign sigmoid_table_675_7_sva_dfm_1 = sigmoid_table_675_7_sva | (~ initialized_sva);
  assign sigmoid_table_676_7_sva_dfm_1 = sigmoid_table_676_7_sva | (~ initialized_sva);
  assign sigmoid_table_677_7_sva_dfm_1 = sigmoid_table_677_7_sva | (~ initialized_sva);
  assign sigmoid_table_678_7_sva_dfm_1 = sigmoid_table_678_7_sva | (~ initialized_sva);
  assign sigmoid_table_679_7_sva_dfm_1 = sigmoid_table_679_7_sva | (~ initialized_sva);
  assign sigmoid_table_680_7_sva_dfm_1 = sigmoid_table_680_7_sva | (~ initialized_sva);
  assign sigmoid_table_681_7_sva_dfm_1 = sigmoid_table_681_7_sva | (~ initialized_sva);
  assign sigmoid_table_682_7_sva_dfm_1 = sigmoid_table_682_7_sva | (~ initialized_sva);
  assign sigmoid_table_683_7_sva_dfm_1 = sigmoid_table_683_7_sva | (~ initialized_sva);
  assign sigmoid_table_684_7_sva_dfm_1 = sigmoid_table_684_7_sva | (~ initialized_sva);
  assign sigmoid_table_685_7_sva_dfm_1 = sigmoid_table_685_7_sva | (~ initialized_sva);
  assign sigmoid_table_686_6_sva_dfm_1 = sigmoid_table_686_6_sva | (~ initialized_sva);
  assign sigmoid_table_687_6_sva_dfm_1 = sigmoid_table_687_6_sva | (~ initialized_sva);
  assign sigmoid_table_688_6_sva_dfm_1 = sigmoid_table_688_6_sva | (~ initialized_sva);
  assign sigmoid_table_689_6_sva_dfm_1 = sigmoid_table_689_6_sva | (~ initialized_sva);
  assign sigmoid_table_690_6_sva_dfm_1 = sigmoid_table_690_6_sva | (~ initialized_sva);
  assign sigmoid_table_691_6_sva_dfm_1 = sigmoid_table_691_6_sva | (~ initialized_sva);
  assign sigmoid_table_692_6_sva_dfm_1 = sigmoid_table_692_6_sva | (~ initialized_sva);
  assign sigmoid_table_693_6_sva_dfm_1 = sigmoid_table_693_6_sva | (~ initialized_sva);
  assign sigmoid_table_694_6_sva_dfm_1 = sigmoid_table_694_6_sva | (~ initialized_sva);
  assign sigmoid_table_695_6_sva_dfm_1 = sigmoid_table_695_6_sva | (~ initialized_sva);
  assign sigmoid_table_696_6_sva_dfm_1 = sigmoid_table_696_6_sva | (~ initialized_sva);
  assign sigmoid_table_697_6_sva_dfm_1 = sigmoid_table_697_6_sva | (~ initialized_sva);
  assign sigmoid_table_698_6_sva_dfm_1 = sigmoid_table_698_6_sva | (~ initialized_sva);
  assign sigmoid_table_699_6_sva_dfm_1 = sigmoid_table_699_6_sva | (~ initialized_sva);
  assign sigmoid_table_700_6_sva_dfm_1 = sigmoid_table_700_6_sva | (~ initialized_sva);
  assign sigmoid_table_701_6_sva_dfm_1 = sigmoid_table_701_6_sva | (~ initialized_sva);
  assign sigmoid_table_702_6_sva_dfm_1 = sigmoid_table_702_6_sva | (~ initialized_sva);
  assign sigmoid_table_703_6_sva_dfm_1 = sigmoid_table_703_6_sva | (~ initialized_sva);
  assign sigmoid_table_704_6_sva_dfm_1 = sigmoid_table_704_6_sva | (~ initialized_sva);
  assign sigmoid_table_705_6_sva_dfm_1 = sigmoid_table_705_6_sva | (~ initialized_sva);
  assign sigmoid_table_706_6_sva_dfm_1 = sigmoid_table_706_6_sva | (~ initialized_sva);
  assign sigmoid_table_707_6_sva_dfm_1 = sigmoid_table_707_6_sva | (~ initialized_sva);
  assign sigmoid_table_708_6_sva_dfm_1 = sigmoid_table_708_6_sva | (~ initialized_sva);
  assign sigmoid_table_709_6_sva_dfm_1 = sigmoid_table_709_6_sva | (~ initialized_sva);
  assign sigmoid_table_710_6_sva_dfm_1 = sigmoid_table_710_6_sva | (~ initialized_sva);
  assign sigmoid_table_711_6_sva_dfm_1 = sigmoid_table_711_6_sva | (~ initialized_sva);
  assign sigmoid_table_712_6_sva_dfm_1 = sigmoid_table_712_6_sva | (~ initialized_sva);
  assign sigmoid_table_713_6_sva_dfm_1 = sigmoid_table_713_6_sva | (~ initialized_sva);
  assign sigmoid_table_714_6_sva_dfm_1 = sigmoid_table_714_6_sva | (~ initialized_sva);
  assign sigmoid_table_715_6_sva_dfm_1 = sigmoid_table_715_6_sva | (~ initialized_sva);
  assign sigmoid_table_716_6_sva_dfm_1 = sigmoid_table_716_6_sva | (~ initialized_sva);
  assign sigmoid_table_717_6_sva_dfm_1 = sigmoid_table_717_6_sva | (~ initialized_sva);
  assign sigmoid_table_718_6_sva_dfm_1 = sigmoid_table_718_6_sva | (~ initialized_sva);
  assign sigmoid_table_719_6_sva_dfm_1 = sigmoid_table_719_6_sva | (~ initialized_sva);
  assign sigmoid_table_720_6_sva_dfm_1 = sigmoid_table_720_6_sva | (~ initialized_sva);
  assign sigmoid_table_721_6_sva_dfm_1 = sigmoid_table_721_6_sva | (~ initialized_sva);
  assign sigmoid_table_722_6_sva_dfm_1 = sigmoid_table_722_6_sva | (~ initialized_sva);
  assign sigmoid_table_723_6_sva_dfm_1 = sigmoid_table_723_6_sva | (~ initialized_sva);
  assign sigmoid_table_724_6_sva_dfm_1 = sigmoid_table_724_6_sva | (~ initialized_sva);
  assign sigmoid_table_725_6_sva_dfm_1 = sigmoid_table_725_6_sva | (~ initialized_sva);
  assign sigmoid_table_726_6_sva_dfm_1 = sigmoid_table_726_6_sva | (~ initialized_sva);
  assign sigmoid_table_727_6_sva_dfm_1 = sigmoid_table_727_6_sva | (~ initialized_sva);
  assign sigmoid_table_728_6_sva_dfm_1 = sigmoid_table_728_6_sva | (~ initialized_sva);
  assign sigmoid_table_729_6_sva_dfm_1 = sigmoid_table_729_6_sva | (~ initialized_sva);
  assign sigmoid_table_730_6_sva_dfm_1 = sigmoid_table_730_6_sva | (~ initialized_sva);
  assign sigmoid_table_731_6_sva_dfm_1 = sigmoid_table_731_6_sva | (~ initialized_sva);
  assign sigmoid_table_732_5_sva_dfm_1 = sigmoid_table_732_5_sva | (~ initialized_sva);
  assign sigmoid_table_733_5_sva_dfm_1 = sigmoid_table_733_5_sva | (~ initialized_sva);
  assign sigmoid_table_734_5_sva_dfm_1 = sigmoid_table_734_5_sva | (~ initialized_sva);
  assign sigmoid_table_735_5_sva_dfm_1 = sigmoid_table_735_5_sva | (~ initialized_sva);
  assign sigmoid_table_736_5_sva_dfm_1 = sigmoid_table_736_5_sva | (~ initialized_sva);
  assign sigmoid_table_737_5_sva_dfm_1 = sigmoid_table_737_5_sva | (~ initialized_sva);
  assign sigmoid_table_738_5_sva_dfm_1 = sigmoid_table_738_5_sva | (~ initialized_sva);
  assign sigmoid_table_739_5_sva_dfm_1 = sigmoid_table_739_5_sva | (~ initialized_sva);
  assign sigmoid_table_740_5_sva_dfm_1 = sigmoid_table_740_5_sva | (~ initialized_sva);
  assign sigmoid_table_741_5_sva_dfm_1 = sigmoid_table_741_5_sva | (~ initialized_sva);
  assign sigmoid_table_742_5_sva_dfm_1 = sigmoid_table_742_5_sva | (~ initialized_sva);
  assign sigmoid_table_743_5_sva_dfm_1 = sigmoid_table_743_5_sva | (~ initialized_sva);
  assign sigmoid_table_744_5_sva_dfm_1 = sigmoid_table_744_5_sva | (~ initialized_sva);
  assign sigmoid_table_745_5_sva_dfm_1 = sigmoid_table_745_5_sva | (~ initialized_sva);
  assign sigmoid_table_746_5_sva_dfm_1 = sigmoid_table_746_5_sva | (~ initialized_sva);
  assign sigmoid_table_747_5_sva_dfm_1 = sigmoid_table_747_5_sva | (~ initialized_sva);
  assign sigmoid_table_748_5_sva_dfm_1 = sigmoid_table_748_5_sva | (~ initialized_sva);
  assign sigmoid_table_749_5_sva_dfm_1 = sigmoid_table_749_5_sva | (~ initialized_sva);
  assign sigmoid_table_750_5_sva_dfm_1 = sigmoid_table_750_5_sva | (~ initialized_sva);
  assign sigmoid_table_751_5_sva_dfm_1 = sigmoid_table_751_5_sva | (~ initialized_sva);
  assign sigmoid_table_752_5_sva_dfm_1 = sigmoid_table_752_5_sva | (~ initialized_sva);
  assign sigmoid_table_753_5_sva_dfm_1 = sigmoid_table_753_5_sva | (~ initialized_sva);
  assign sigmoid_table_754_5_sva_dfm_1 = sigmoid_table_754_5_sva | (~ initialized_sva);
  assign sigmoid_table_755_5_sva_dfm_1 = sigmoid_table_755_5_sva | (~ initialized_sva);
  assign sigmoid_table_756_5_sva_dfm_1 = sigmoid_table_756_5_sva | (~ initialized_sva);
  assign sigmoid_table_757_5_sva_dfm_1 = sigmoid_table_757_5_sva | (~ initialized_sva);
  assign sigmoid_table_758_5_sva_dfm_1 = sigmoid_table_758_5_sva | (~ initialized_sva);
  assign sigmoid_table_759_5_sva_dfm_1 = sigmoid_table_759_5_sva | (~ initialized_sva);
  assign sigmoid_table_760_5_sva_dfm_1 = sigmoid_table_760_5_sva | (~ initialized_sva);
  assign sigmoid_table_761_5_sva_dfm_1 = sigmoid_table_761_5_sva | (~ initialized_sva);
  assign sigmoid_table_762_5_sva_dfm_1 = sigmoid_table_762_5_sva | (~ initialized_sva);
  assign sigmoid_table_763_5_sva_dfm_1 = sigmoid_table_763_5_sva | (~ initialized_sva);
  assign sigmoid_table_764_5_sva_dfm_1 = sigmoid_table_764_5_sva | (~ initialized_sva);
  assign sigmoid_table_765_5_sva_dfm_1 = sigmoid_table_765_5_sva | (~ initialized_sva);
  assign sigmoid_table_766_5_sva_dfm_1 = sigmoid_table_766_5_sva | (~ initialized_sva);
  assign sigmoid_table_767_5_sva_dfm_1 = sigmoid_table_767_5_sva | (~ initialized_sva);
  assign sigmoid_table_768_5_sva_dfm_1 = sigmoid_table_768_5_sva | (~ initialized_sva);
  assign sigmoid_table_769_5_sva_dfm_1 = sigmoid_table_769_5_sva | (~ initialized_sva);
  assign sigmoid_table_770_5_sva_dfm_1 = sigmoid_table_770_5_sva | (~ initialized_sva);
  assign sigmoid_table_771_5_sva_dfm_1 = sigmoid_table_771_5_sva | (~ initialized_sva);
  assign sigmoid_table_772_5_sva_dfm_1 = sigmoid_table_772_5_sva | (~ initialized_sva);
  assign sigmoid_table_773_5_sva_dfm_1 = sigmoid_table_773_5_sva | (~ initialized_sva);
  assign sigmoid_table_774_5_sva_dfm_1 = sigmoid_table_774_5_sva | (~ initialized_sva);
  assign sigmoid_table_775_5_sva_dfm_1 = sigmoid_table_775_5_sva | (~ initialized_sva);
  assign sigmoid_table_776_5_sva_dfm_1 = sigmoid_table_776_5_sva | (~ initialized_sva);
  assign sigmoid_table_777_5_sva_dfm_1 = sigmoid_table_777_5_sva | (~ initialized_sva);
  assign sigmoid_table_778_4_sva_dfm_1 = sigmoid_table_778_4_sva | (~ initialized_sva);
  assign sigmoid_table_779_4_sva_dfm_1 = sigmoid_table_779_4_sva | (~ initialized_sva);
  assign sigmoid_table_780_4_sva_dfm_1 = sigmoid_table_780_4_sva | (~ initialized_sva);
  assign sigmoid_table_781_4_sva_dfm_1 = sigmoid_table_781_4_sva | (~ initialized_sva);
  assign sigmoid_table_782_4_sva_dfm_1 = sigmoid_table_782_4_sva | (~ initialized_sva);
  assign sigmoid_table_783_4_sva_dfm_1 = sigmoid_table_783_4_sva | (~ initialized_sva);
  assign sigmoid_table_784_4_sva_dfm_1 = sigmoid_table_784_4_sva | (~ initialized_sva);
  assign sigmoid_table_785_4_sva_dfm_1 = sigmoid_table_785_4_sva | (~ initialized_sva);
  assign sigmoid_table_786_4_sva_dfm_1 = sigmoid_table_786_4_sva | (~ initialized_sva);
  assign sigmoid_table_787_4_sva_dfm_1 = sigmoid_table_787_4_sva | (~ initialized_sva);
  assign sigmoid_table_788_4_sva_dfm_1 = sigmoid_table_788_4_sva | (~ initialized_sva);
  assign sigmoid_table_789_4_sva_dfm_1 = sigmoid_table_789_4_sva | (~ initialized_sva);
  assign sigmoid_table_790_4_sva_dfm_1 = sigmoid_table_790_4_sva | (~ initialized_sva);
  assign sigmoid_table_791_4_sva_dfm_1 = sigmoid_table_791_4_sva | (~ initialized_sva);
  assign sigmoid_table_792_4_sva_dfm_1 = sigmoid_table_792_4_sva | (~ initialized_sva);
  assign sigmoid_table_793_4_sva_dfm_1 = sigmoid_table_793_4_sva | (~ initialized_sva);
  assign sigmoid_table_794_4_sva_dfm_1 = sigmoid_table_794_4_sva | (~ initialized_sva);
  assign sigmoid_table_795_4_sva_dfm_1 = sigmoid_table_795_4_sva | (~ initialized_sva);
  assign sigmoid_table_796_4_sva_dfm_1 = sigmoid_table_796_4_sva | (~ initialized_sva);
  assign sigmoid_table_797_4_sva_dfm_1 = sigmoid_table_797_4_sva | (~ initialized_sva);
  assign sigmoid_table_798_4_sva_dfm_1 = sigmoid_table_798_4_sva | (~ initialized_sva);
  assign sigmoid_table_799_4_sva_dfm_1 = sigmoid_table_799_4_sva | (~ initialized_sva);
  assign sigmoid_table_800_4_sva_dfm_1 = sigmoid_table_800_4_sva | (~ initialized_sva);
  assign sigmoid_table_801_4_sva_dfm_1 = sigmoid_table_801_4_sva | (~ initialized_sva);
  assign sigmoid_table_802_4_sva_dfm_1 = sigmoid_table_802_4_sva | (~ initialized_sva);
  assign sigmoid_table_803_4_sva_dfm_1 = sigmoid_table_803_4_sva | (~ initialized_sva);
  assign sigmoid_table_804_4_sva_dfm_1 = sigmoid_table_804_4_sva | (~ initialized_sva);
  assign sigmoid_table_805_4_sva_dfm_1 = sigmoid_table_805_4_sva | (~ initialized_sva);
  assign sigmoid_table_806_4_sva_dfm_1 = sigmoid_table_806_4_sva | (~ initialized_sva);
  assign sigmoid_table_807_4_sva_dfm_1 = sigmoid_table_807_4_sva | (~ initialized_sva);
  assign sigmoid_table_808_4_sva_dfm_1 = sigmoid_table_808_4_sva | (~ initialized_sva);
  assign sigmoid_table_809_4_sva_dfm_1 = sigmoid_table_809_4_sva | (~ initialized_sva);
  assign sigmoid_table_810_4_sva_dfm_1 = sigmoid_table_810_4_sva | (~ initialized_sva);
  assign sigmoid_table_811_4_sva_dfm_1 = sigmoid_table_811_4_sva | (~ initialized_sva);
  assign sigmoid_table_812_4_sva_dfm_1 = sigmoid_table_812_4_sva | (~ initialized_sva);
  assign sigmoid_table_813_4_sva_dfm_1 = sigmoid_table_813_4_sva | (~ initialized_sva);
  assign sigmoid_table_814_4_sva_dfm_1 = sigmoid_table_814_4_sva | (~ initialized_sva);
  assign sigmoid_table_815_4_sva_dfm_1 = sigmoid_table_815_4_sva | (~ initialized_sva);
  assign sigmoid_table_816_4_sva_dfm_1 = sigmoid_table_816_4_sva | (~ initialized_sva);
  assign sigmoid_table_817_4_sva_dfm_1 = sigmoid_table_817_4_sva | (~ initialized_sva);
  assign sigmoid_table_818_4_sva_dfm_1 = sigmoid_table_818_4_sva | (~ initialized_sva);
  assign sigmoid_table_819_4_sva_dfm_1 = sigmoid_table_819_4_sva | (~ initialized_sva);
  assign sigmoid_table_820_4_sva_dfm_1 = sigmoid_table_820_4_sva | (~ initialized_sva);
  assign sigmoid_table_821_4_sva_dfm_1 = sigmoid_table_821_4_sva | (~ initialized_sva);
  assign sigmoid_table_822_3_sva_dfm_1 = sigmoid_table_822_3_sva | (~ initialized_sva);
  assign sigmoid_table_823_3_sva_dfm_1 = sigmoid_table_823_3_sva | (~ initialized_sva);
  assign sigmoid_table_824_3_sva_dfm_1 = sigmoid_table_824_3_sva | (~ initialized_sva);
  assign sigmoid_table_825_3_sva_dfm_1 = sigmoid_table_825_3_sva | (~ initialized_sva);
  assign sigmoid_table_826_3_sva_dfm_1 = sigmoid_table_826_3_sva | (~ initialized_sva);
  assign sigmoid_table_827_3_sva_dfm_1 = sigmoid_table_827_3_sva | (~ initialized_sva);
  assign sigmoid_table_828_3_sva_dfm_1 = sigmoid_table_828_3_sva | (~ initialized_sva);
  assign sigmoid_table_829_3_sva_dfm_1 = sigmoid_table_829_3_sva | (~ initialized_sva);
  assign sigmoid_table_830_3_sva_dfm_1 = sigmoid_table_830_3_sva | (~ initialized_sva);
  assign sigmoid_table_831_3_sva_dfm_1 = sigmoid_table_831_3_sva | (~ initialized_sva);
  assign sigmoid_table_832_3_sva_dfm_1 = sigmoid_table_832_3_sva | (~ initialized_sva);
  assign sigmoid_table_833_3_sva_dfm_1 = sigmoid_table_833_3_sva | (~ initialized_sva);
  assign sigmoid_table_834_3_sva_dfm_1 = sigmoid_table_834_3_sva | (~ initialized_sva);
  assign sigmoid_table_835_3_sva_dfm_1 = sigmoid_table_835_3_sva | (~ initialized_sva);
  assign sigmoid_table_836_3_sva_dfm_1 = sigmoid_table_836_3_sva | (~ initialized_sva);
  assign sigmoid_table_837_3_sva_dfm_1 = sigmoid_table_837_3_sva | (~ initialized_sva);
  assign sigmoid_table_838_3_sva_dfm_1 = sigmoid_table_838_3_sva | (~ initialized_sva);
  assign sigmoid_table_839_3_sva_dfm_1 = sigmoid_table_839_3_sva | (~ initialized_sva);
  assign sigmoid_table_840_3_sva_dfm_1 = sigmoid_table_840_3_sva | (~ initialized_sva);
  assign sigmoid_table_841_3_sva_dfm_1 = sigmoid_table_841_3_sva | (~ initialized_sva);
  assign sigmoid_table_842_3_sva_dfm_1 = sigmoid_table_842_3_sva | (~ initialized_sva);
  assign sigmoid_table_843_3_sva_dfm_1 = sigmoid_table_843_3_sva | (~ initialized_sva);
  assign sigmoid_table_844_3_sva_dfm_1 = sigmoid_table_844_3_sva | (~ initialized_sva);
  assign sigmoid_table_845_3_sva_dfm_1 = sigmoid_table_845_3_sva | (~ initialized_sva);
  assign sigmoid_table_846_3_sva_dfm_1 = sigmoid_table_846_3_sva | (~ initialized_sva);
  assign sigmoid_table_847_3_sva_dfm_1 = sigmoid_table_847_3_sva | (~ initialized_sva);
  assign sigmoid_table_848_3_sva_dfm_1 = sigmoid_table_848_3_sva | (~ initialized_sva);
  assign sigmoid_table_849_3_sva_dfm_1 = sigmoid_table_849_3_sva | (~ initialized_sva);
  assign sigmoid_table_850_3_sva_dfm_1 = sigmoid_table_850_3_sva | (~ initialized_sva);
  assign sigmoid_table_851_3_sva_dfm_1 = sigmoid_table_851_3_sva | (~ initialized_sva);
  assign sigmoid_table_852_3_sva_dfm_1 = sigmoid_table_852_3_sva | (~ initialized_sva);
  assign sigmoid_table_853_3_sva_dfm_1 = sigmoid_table_853_3_sva | (~ initialized_sva);
  assign sigmoid_table_854_3_sva_dfm_1 = sigmoid_table_854_3_sva | (~ initialized_sva);
  assign sigmoid_table_855_3_sva_dfm_1 = sigmoid_table_855_3_sva | (~ initialized_sva);
  assign sigmoid_table_856_3_sva_dfm_1 = sigmoid_table_856_3_sva | (~ initialized_sva);
  assign sigmoid_table_857_3_sva_dfm_1 = sigmoid_table_857_3_sva | (~ initialized_sva);
  assign sigmoid_table_858_3_sva_dfm_1 = sigmoid_table_858_3_sva | (~ initialized_sva);
  assign sigmoid_table_859_3_sva_dfm_1 = sigmoid_table_859_3_sva | (~ initialized_sva);
  assign sigmoid_table_860_3_sva_dfm_1 = sigmoid_table_860_3_sva | (~ initialized_sva);
  assign sigmoid_table_861_3_sva_dfm_1 = sigmoid_table_861_3_sva | (~ initialized_sva);
  assign sigmoid_table_862_3_sva_dfm_1 = sigmoid_table_862_3_sva | (~ initialized_sva);
  assign sigmoid_table_863_3_sva_dfm_1 = sigmoid_table_863_3_sva | (~ initialized_sva);
  assign sigmoid_table_864_3_sva_dfm_1 = sigmoid_table_864_3_sva | (~ initialized_sva);
  assign sigmoid_table_865_3_sva_dfm_1 = sigmoid_table_865_3_sva | (~ initialized_sva);
  assign sigmoid_table_866_3_sva_dfm_1 = sigmoid_table_866_3_sva | (~ initialized_sva);
  assign sigmoid_table_867_2_sva_dfm_1 = sigmoid_table_867_2_sva | (~ initialized_sva);
  assign sigmoid_table_868_2_sva_dfm_1 = sigmoid_table_868_2_sva | (~ initialized_sva);
  assign sigmoid_table_869_2_sva_dfm_1 = sigmoid_table_869_2_sva | (~ initialized_sva);
  assign sigmoid_table_870_2_sva_dfm_1 = sigmoid_table_870_2_sva | (~ initialized_sva);
  assign sigmoid_table_871_2_sva_dfm_1 = sigmoid_table_871_2_sva | (~ initialized_sva);
  assign sigmoid_table_872_2_sva_dfm_1 = sigmoid_table_872_2_sva | (~ initialized_sva);
  assign sigmoid_table_873_2_sva_dfm_1 = sigmoid_table_873_2_sva | (~ initialized_sva);
  assign sigmoid_table_874_2_sva_dfm_1 = sigmoid_table_874_2_sva | (~ initialized_sva);
  assign sigmoid_table_875_2_sva_dfm_1 = sigmoid_table_875_2_sva | (~ initialized_sva);
  assign sigmoid_table_876_2_sva_dfm_1 = sigmoid_table_876_2_sva | (~ initialized_sva);
  assign sigmoid_table_877_2_sva_dfm_1 = sigmoid_table_877_2_sva | (~ initialized_sva);
  assign sigmoid_table_878_2_sva_dfm_1 = sigmoid_table_878_2_sva | (~ initialized_sva);
  assign sigmoid_table_879_2_sva_dfm_1 = sigmoid_table_879_2_sva | (~ initialized_sva);
  assign sigmoid_table_880_2_sva_dfm_1 = sigmoid_table_880_2_sva | (~ initialized_sva);
  assign sigmoid_table_881_2_sva_dfm_1 = sigmoid_table_881_2_sva | (~ initialized_sva);
  assign sigmoid_table_882_2_sva_dfm_1 = sigmoid_table_882_2_sva | (~ initialized_sva);
  assign sigmoid_table_883_2_sva_dfm_1 = sigmoid_table_883_2_sva | (~ initialized_sva);
  assign sigmoid_table_884_2_sva_dfm_1 = sigmoid_table_884_2_sva | (~ initialized_sva);
  assign sigmoid_table_885_2_sva_dfm_1 = sigmoid_table_885_2_sva | (~ initialized_sva);
  assign sigmoid_table_886_2_sva_dfm_1 = sigmoid_table_886_2_sva | (~ initialized_sva);
  assign sigmoid_table_887_2_sva_dfm_1 = sigmoid_table_887_2_sva | (~ initialized_sva);
  assign sigmoid_table_888_2_sva_dfm_1 = sigmoid_table_888_2_sva | (~ initialized_sva);
  assign sigmoid_table_889_2_sva_dfm_1 = sigmoid_table_889_2_sva | (~ initialized_sva);
  assign sigmoid_table_890_2_sva_dfm_1 = sigmoid_table_890_2_sva | (~ initialized_sva);
  assign sigmoid_table_891_2_sva_dfm_1 = sigmoid_table_891_2_sva | (~ initialized_sva);
  assign sigmoid_table_892_2_sva_dfm_1 = sigmoid_table_892_2_sva | (~ initialized_sva);
  assign sigmoid_table_893_2_sva_dfm_1 = sigmoid_table_893_2_sva | (~ initialized_sva);
  assign sigmoid_table_894_2_sva_dfm_1 = sigmoid_table_894_2_sva | (~ initialized_sva);
  assign sigmoid_table_895_2_sva_dfm_1 = sigmoid_table_895_2_sva | (~ initialized_sva);
  assign sigmoid_table_896_2_sva_dfm_1 = sigmoid_table_896_2_sva | (~ initialized_sva);
  assign sigmoid_table_897_2_sva_dfm_1 = sigmoid_table_897_2_sva | (~ initialized_sva);
  assign sigmoid_table_898_2_sva_dfm_1 = sigmoid_table_898_2_sva | (~ initialized_sva);
  assign sigmoid_table_899_2_sva_dfm_1 = sigmoid_table_899_2_sva | (~ initialized_sva);
  assign sigmoid_table_900_2_sva_dfm_1 = sigmoid_table_900_2_sva | (~ initialized_sva);
  assign sigmoid_table_901_2_sva_dfm_1 = sigmoid_table_901_2_sva | (~ initialized_sva);
  assign sigmoid_table_902_2_sva_dfm_1 = sigmoid_table_902_2_sva | (~ initialized_sva);
  assign sigmoid_table_903_2_sva_dfm_1 = sigmoid_table_903_2_sva | (~ initialized_sva);
  assign sigmoid_table_904_2_sva_dfm_1 = sigmoid_table_904_2_sva | (~ initialized_sva);
  assign sigmoid_table_905_2_sva_dfm_1 = sigmoid_table_905_2_sva | (~ initialized_sva);
  assign sigmoid_table_906_2_sva_dfm_1 = sigmoid_table_906_2_sva | (~ initialized_sva);
  assign sigmoid_table_907_2_sva_dfm_1 = sigmoid_table_907_2_sva | (~ initialized_sva);
  assign sigmoid_table_908_2_sva_dfm_1 = sigmoid_table_908_2_sva | (~ initialized_sva);
  assign sigmoid_table_909_2_sva_dfm_1 = sigmoid_table_909_2_sva | (~ initialized_sva);
  assign sigmoid_table_910_2_sva_dfm_1 = sigmoid_table_910_2_sva | (~ initialized_sva);
  assign sigmoid_table_911_1_sva_dfm_1 = sigmoid_table_911_1_sva | (~ initialized_sva);
  assign sigmoid_table_912_1_sva_dfm_1 = sigmoid_table_912_1_sva | (~ initialized_sva);
  assign sigmoid_table_913_1_sva_dfm_1 = sigmoid_table_913_1_sva | (~ initialized_sva);
  assign sigmoid_table_914_1_sva_dfm_1 = sigmoid_table_914_1_sva | (~ initialized_sva);
  assign sigmoid_table_915_1_sva_dfm_1 = sigmoid_table_915_1_sva | (~ initialized_sva);
  assign sigmoid_table_916_1_sva_dfm_1 = sigmoid_table_916_1_sva | (~ initialized_sva);
  assign sigmoid_table_917_1_sva_dfm_1 = sigmoid_table_917_1_sva | (~ initialized_sva);
  assign sigmoid_table_918_1_sva_dfm_1 = sigmoid_table_918_1_sva | (~ initialized_sva);
  assign sigmoid_table_919_1_sva_dfm_1 = sigmoid_table_919_1_sva | (~ initialized_sva);
  assign sigmoid_table_920_1_sva_dfm_1 = sigmoid_table_920_1_sva | (~ initialized_sva);
  assign sigmoid_table_921_1_sva_dfm_1 = sigmoid_table_921_1_sva | (~ initialized_sva);
  assign sigmoid_table_922_1_sva_dfm_1 = sigmoid_table_922_1_sva | (~ initialized_sva);
  assign sigmoid_table_923_1_sva_dfm_1 = sigmoid_table_923_1_sva | (~ initialized_sva);
  assign sigmoid_table_924_1_sva_dfm_1 = sigmoid_table_924_1_sva | (~ initialized_sva);
  assign sigmoid_table_925_1_sva_dfm_1 = sigmoid_table_925_1_sva | (~ initialized_sva);
  assign sigmoid_table_926_1_sva_dfm_1 = sigmoid_table_926_1_sva | (~ initialized_sva);
  assign sigmoid_table_927_1_sva_dfm_1 = sigmoid_table_927_1_sva | (~ initialized_sva);
  assign sigmoid_table_928_1_sva_dfm_1 = sigmoid_table_928_1_sva | (~ initialized_sva);
  assign sigmoid_table_929_1_sva_dfm_1 = sigmoid_table_929_1_sva | (~ initialized_sva);
  assign sigmoid_table_930_1_sva_dfm_1 = sigmoid_table_930_1_sva | (~ initialized_sva);
  assign sigmoid_table_931_1_sva_dfm_1 = sigmoid_table_931_1_sva | (~ initialized_sva);
  assign sigmoid_table_932_1_sva_dfm_1 = sigmoid_table_932_1_sva | (~ initialized_sva);
  assign sigmoid_table_933_1_sva_dfm_1 = sigmoid_table_933_1_sva | (~ initialized_sva);
  assign sigmoid_table_934_1_sva_dfm_1 = sigmoid_table_934_1_sva | (~ initialized_sva);
  assign sigmoid_table_935_1_sva_dfm_1 = sigmoid_table_935_1_sva | (~ initialized_sva);
  assign sigmoid_table_936_1_sva_dfm_1 = sigmoid_table_936_1_sva | (~ initialized_sva);
  assign sigmoid_table_937_1_sva_dfm_1 = sigmoid_table_937_1_sva | (~ initialized_sva);
  assign sigmoid_table_938_1_sva_dfm_1 = sigmoid_table_938_1_sva | (~ initialized_sva);
  assign sigmoid_table_939_1_sva_dfm_1 = sigmoid_table_939_1_sva | (~ initialized_sva);
  assign sigmoid_table_940_1_sva_dfm_1 = sigmoid_table_940_1_sva | (~ initialized_sva);
  assign sigmoid_table_941_1_sva_dfm_1 = sigmoid_table_941_1_sva | (~ initialized_sva);
  assign sigmoid_table_942_1_sva_dfm_1 = sigmoid_table_942_1_sva | (~ initialized_sva);
  assign sigmoid_table_943_1_sva_dfm_1 = sigmoid_table_943_1_sva | (~ initialized_sva);
  assign sigmoid_table_944_1_sva_dfm_1 = sigmoid_table_944_1_sva | (~ initialized_sva);
  assign sigmoid_table_945_1_sva_dfm_1 = sigmoid_table_945_1_sva | (~ initialized_sva);
  assign sigmoid_table_946_1_sva_dfm_1 = sigmoid_table_946_1_sva | (~ initialized_sva);
  assign sigmoid_table_947_1_sva_dfm_1 = sigmoid_table_947_1_sva | (~ initialized_sva);
  assign sigmoid_table_948_1_sva_dfm_1 = sigmoid_table_948_1_sva | (~ initialized_sva);
  assign sigmoid_table_949_1_sva_dfm_1 = sigmoid_table_949_1_sva | (~ initialized_sva);
  assign sigmoid_table_950_1_sva_dfm_1 = sigmoid_table_950_1_sva | (~ initialized_sva);
  assign sigmoid_table_951_1_sva_dfm_1 = sigmoid_table_951_1_sva | (~ initialized_sva);
  assign sigmoid_table_952_1_sva_dfm_1 = sigmoid_table_952_1_sva | (~ initialized_sva);
  assign sigmoid_table_953_1_sva_dfm_1 = sigmoid_table_953_1_sva | (~ initialized_sva);
  assign sigmoid_table_954_1_sva_dfm_1 = sigmoid_table_954_1_sva | (~ initialized_sva);
  assign sigmoid_table_113_1_sva_dfm_1 = sigmoid_table_113_1_sva | (~ initialized_sva);
  assign sigmoid_table_114_1_sva_dfm_1 = sigmoid_table_114_1_sva | (~ initialized_sva);
  assign sigmoid_table_115_1_sva_dfm_1 = sigmoid_table_115_1_sva | (~ initialized_sva);
  assign sigmoid_table_116_1_sva_dfm_1 = sigmoid_table_116_1_sva | (~ initialized_sva);
  assign sigmoid_table_117_1_sva_dfm_1 = sigmoid_table_117_1_sva | (~ initialized_sva);
  assign sigmoid_table_118_1_sva_dfm_1 = sigmoid_table_118_1_sva | (~ initialized_sva);
  assign sigmoid_table_119_1_sva_dfm_1 = sigmoid_table_119_1_sva | (~ initialized_sva);
  assign sigmoid_table_120_1_sva_dfm_1 = sigmoid_table_120_1_sva | (~ initialized_sva);
  assign sigmoid_table_121_1_sva_dfm_1 = sigmoid_table_121_1_sva | (~ initialized_sva);
  assign sigmoid_table_122_1_sva_dfm_1 = sigmoid_table_122_1_sva | (~ initialized_sva);
  assign sigmoid_table_123_1_sva_dfm_1 = sigmoid_table_123_1_sva | (~ initialized_sva);
  assign sigmoid_table_124_1_sva_dfm_1 = sigmoid_table_124_1_sva | (~ initialized_sva);
  assign sigmoid_table_125_1_sva_dfm_1 = sigmoid_table_125_1_sva | (~ initialized_sva);
  assign sigmoid_table_126_1_sva_dfm_1 = sigmoid_table_126_1_sva | (~ initialized_sva);
  assign sigmoid_table_127_1_sva_dfm_1 = sigmoid_table_127_1_sva | (~ initialized_sva);
  assign sigmoid_table_128_1_sva_dfm_1 = sigmoid_table_128_1_sva | (~ initialized_sva);
  assign sigmoid_table_129_1_sva_dfm_1 = sigmoid_table_129_1_sva | (~ initialized_sva);
  assign sigmoid_table_130_1_sva_dfm_1 = sigmoid_table_130_1_sva | (~ initialized_sva);
  assign sigmoid_table_131_1_sva_dfm_1 = sigmoid_table_131_1_sva | (~ initialized_sva);
  assign sigmoid_table_132_1_sva_dfm_1 = sigmoid_table_132_1_sva | (~ initialized_sva);
  assign sigmoid_table_133_1_sva_dfm_1 = sigmoid_table_133_1_sva | (~ initialized_sva);
  assign sigmoid_table_134_1_sva_dfm_1 = sigmoid_table_134_1_sva | (~ initialized_sva);
  assign sigmoid_table_135_1_sva_dfm_1 = sigmoid_table_135_1_sva | (~ initialized_sva);
  assign sigmoid_table_136_1_sva_dfm_1 = sigmoid_table_136_1_sva | (~ initialized_sva);
  assign sigmoid_table_137_1_sva_dfm_1 = sigmoid_table_137_1_sva | (~ initialized_sva);
  assign sigmoid_table_138_1_sva_dfm_1 = sigmoid_table_138_1_sva | (~ initialized_sva);
  assign sigmoid_table_184_1_sva_dfm_1 = sigmoid_table_184_1_sva | (~ initialized_sva);
  assign sigmoid_table_185_1_sva_dfm_1 = sigmoid_table_185_1_sva | (~ initialized_sva);
  assign sigmoid_table_186_1_sva_dfm_1 = sigmoid_table_186_1_sva | (~ initialized_sva);
  assign sigmoid_table_187_1_sva_dfm_1 = sigmoid_table_187_1_sva | (~ initialized_sva);
  assign sigmoid_table_188_1_sva_dfm_1 = sigmoid_table_188_1_sva | (~ initialized_sva);
  assign sigmoid_table_189_1_sva_dfm_1 = sigmoid_table_189_1_sva | (~ initialized_sva);
  assign sigmoid_table_190_1_sva_dfm_1 = sigmoid_table_190_1_sva | (~ initialized_sva);
  assign sigmoid_table_191_1_sva_dfm_1 = sigmoid_table_191_1_sva | (~ initialized_sva);
  assign sigmoid_table_192_1_sva_dfm_1 = sigmoid_table_192_1_sva | (~ initialized_sva);
  assign sigmoid_table_193_1_sva_dfm_1 = sigmoid_table_193_1_sva | (~ initialized_sva);
  assign sigmoid_table_217_1_sva_dfm_1 = sigmoid_table_217_1_sva | (~ initialized_sva);
  assign sigmoid_table_218_1_sva_dfm_1 = sigmoid_table_218_1_sva | (~ initialized_sva);
  assign sigmoid_table_219_1_sva_dfm_1 = sigmoid_table_219_1_sva | (~ initialized_sva);
  assign sigmoid_table_220_1_sva_dfm_1 = sigmoid_table_220_1_sva | (~ initialized_sva);
  assign sigmoid_table_221_1_sva_dfm_1 = sigmoid_table_221_1_sva | (~ initialized_sva);
  assign sigmoid_table_222_1_sva_dfm_1 = sigmoid_table_222_1_sva | (~ initialized_sva);
  assign sigmoid_table_239_1_sva_dfm_1 = sigmoid_table_239_1_sva | (~ initialized_sva);
  assign sigmoid_table_240_1_sva_dfm_1 = sigmoid_table_240_1_sva | (~ initialized_sva);
  assign sigmoid_table_241_1_sva_dfm_1 = sigmoid_table_241_1_sva | (~ initialized_sva);
  assign sigmoid_table_242_1_sva_dfm_1 = sigmoid_table_242_1_sva | (~ initialized_sva);
  assign sigmoid_table_255_1_sva_dfm_1 = sigmoid_table_255_1_sva | (~ initialized_sva);
  assign sigmoid_table_256_1_sva_dfm_1 = sigmoid_table_256_1_sva | (~ initialized_sva);
  assign sigmoid_table_257_1_sva_dfm_1 = sigmoid_table_257_1_sva | (~ initialized_sva);
  assign sigmoid_table_258_1_sva_dfm_1 = sigmoid_table_258_1_sva | (~ initialized_sva);
  assign sigmoid_table_268_1_sva_dfm_1 = sigmoid_table_268_1_sva | (~ initialized_sva);
  assign sigmoid_table_269_1_sva_dfm_1 = sigmoid_table_269_1_sva | (~ initialized_sva);
  assign sigmoid_table_270_1_sva_dfm_1 = sigmoid_table_270_1_sva | (~ initialized_sva);
  assign sigmoid_table_279_1_sva_dfm_1 = sigmoid_table_279_1_sva | (~ initialized_sva);
  assign sigmoid_table_280_1_sva_dfm_1 = sigmoid_table_280_1_sva | (~ initialized_sva);
  assign sigmoid_table_281_1_sva_dfm_1 = sigmoid_table_281_1_sva | (~ initialized_sva);
  assign sigmoid_table_288_1_sva_dfm_1 = sigmoid_table_288_1_sva | (~ initialized_sva);
  assign sigmoid_table_289_1_sva_dfm_1 = sigmoid_table_289_1_sva | (~ initialized_sva);
  assign sigmoid_table_290_1_sva_dfm_1 = sigmoid_table_290_1_sva | (~ initialized_sva);
  assign sigmoid_table_297_1_sva_dfm_1 = sigmoid_table_297_1_sva | (~ initialized_sva);
  assign sigmoid_table_298_1_sva_dfm_1 = sigmoid_table_298_1_sva | (~ initialized_sva);
  assign sigmoid_table_304_1_sva_dfm_1 = sigmoid_table_304_1_sva | (~ initialized_sva);
  assign sigmoid_table_305_1_sva_dfm_1 = sigmoid_table_305_1_sva | (~ initialized_sva);
  assign sigmoid_table_311_1_sva_dfm_1 = sigmoid_table_311_1_sva | (~ initialized_sva);
  assign sigmoid_table_317_1_sva_dfm_1 = sigmoid_table_317_1_sva | (~ initialized_sva);
  assign sigmoid_table_322_1_sva_dfm_1 = sigmoid_table_322_1_sva | (~ initialized_sva);
  assign sigmoid_table_323_1_sva_dfm_1 = sigmoid_table_323_1_sva | (~ initialized_sva);
  assign sigmoid_table_328_1_sva_dfm_1 = sigmoid_table_328_1_sva | (~ initialized_sva);
  assign sigmoid_table_332_1_sva_dfm_1 = sigmoid_table_332_1_sva | (~ initialized_sva);
  assign sigmoid_table_333_1_sva_dfm_1 = sigmoid_table_333_1_sva | (~ initialized_sva);
  assign sigmoid_table_337_1_sva_dfm_1 = sigmoid_table_337_1_sva | (~ initialized_sva);
  assign sigmoid_table_341_1_sva_dfm_1 = sigmoid_table_341_1_sva | (~ initialized_sva);
  assign sigmoid_table_345_1_sva_dfm_1 = sigmoid_table_345_1_sva | (~ initialized_sva);
  assign sigmoid_table_349_1_sva_dfm_1 = sigmoid_table_349_1_sva | (~ initialized_sva);
  assign sigmoid_table_353_1_sva_dfm_1 = sigmoid_table_353_1_sva | (~ initialized_sva);
  assign sigmoid_table_356_1_sva_dfm_1 = sigmoid_table_356_1_sva | (~ initialized_sva);
  assign sigmoid_table_363_1_sva_dfm_1 = sigmoid_table_363_1_sva | (~ initialized_sva);
  assign sigmoid_table_366_1_sva_dfm_1 = sigmoid_table_366_1_sva | (~ initialized_sva);
  assign sigmoid_table_374_1_sva_dfm_1 = sigmoid_table_374_1_sva | (~ initialized_sva);
  assign sigmoid_table_377_1_sva_dfm_1 = sigmoid_table_377_1_sva | (~ initialized_sva);
  assign sigmoid_table_382_1_sva_dfm_1 = sigmoid_table_382_1_sva | (~ initialized_sva);
  assign sigmoid_table_384_1_sva_dfm_1 = sigmoid_table_384_1_sva | (~ initialized_sva);
  assign sigmoid_table_389_1_sva_dfm_1 = sigmoid_table_389_1_sva | (~ initialized_sva);
  assign sigmoid_table_391_1_sva_dfm_1 = sigmoid_table_391_1_sva | (~ initialized_sva);
  assign sigmoid_table_393_1_sva_dfm_1 = sigmoid_table_393_1_sva | (~ initialized_sva);
  assign sigmoid_table_407_1_sva_dfm_1 = sigmoid_table_407_1_sva | (~ initialized_sva);
  assign sigmoid_table_409_1_sva_dfm_1 = sigmoid_table_409_1_sva | (~ initialized_sva);
  assign sigmoid_table_414_1_sva_dfm_1 = sigmoid_table_414_1_sva | (~ initialized_sva);
  assign sigmoid_table_416_1_sva_dfm_1 = sigmoid_table_416_1_sva | (~ initialized_sva);
  assign sigmoid_table_419_1_sva_dfm_1 = sigmoid_table_419_1_sva | (~ initialized_sva);
  assign sigmoid_table_424_1_sva_dfm_1 = sigmoid_table_424_1_sva | (~ initialized_sva);
  assign sigmoid_table_427_1_sva_dfm_1 = sigmoid_table_427_1_sva | (~ initialized_sva);
  assign sigmoid_table_430_1_sva_dfm_1 = sigmoid_table_430_1_sva | (~ initialized_sva);
  assign sigmoid_table_433_1_sva_dfm_1 = sigmoid_table_433_1_sva | (~ initialized_sva);
  assign sigmoid_table_437_1_sva_dfm_1 = sigmoid_table_437_1_sva | (~ initialized_sva);
  assign sigmoid_table_440_1_sva_dfm_1 = sigmoid_table_440_1_sva | (~ initialized_sva);
  assign sigmoid_table_444_1_sva_dfm_1 = sigmoid_table_444_1_sva | (~ initialized_sva);
  assign sigmoid_table_445_1_sva_dfm_1 = sigmoid_table_445_1_sva | (~ initialized_sva);
  assign sigmoid_table_449_1_sva_dfm_1 = sigmoid_table_449_1_sva | (~ initialized_sva);
  assign sigmoid_table_454_1_sva_dfm_1 = sigmoid_table_454_1_sva | (~ initialized_sva);
  assign sigmoid_table_460_1_sva_dfm_1 = sigmoid_table_460_1_sva | (~ initialized_sva);
  assign sigmoid_table_461_1_sva_dfm_1 = sigmoid_table_461_1_sva | (~ initialized_sva);
  assign sigmoid_table_468_1_sva_dfm_1 = sigmoid_table_468_1_sva | (~ initialized_sva);
  assign sigmoid_table_469_1_sva_dfm_1 = sigmoid_table_469_1_sva | (~ initialized_sva);
  assign sigmoid_table_479_1_sva_dfm_1 = sigmoid_table_479_1_sva | (~ initialized_sva);
  assign sigmoid_table_480_1_sva_dfm_1 = sigmoid_table_480_1_sva | (~ initialized_sva);
  assign sigmoid_table_481_1_sva_dfm_1 = sigmoid_table_481_1_sva | (~ initialized_sva);
  assign sigmoid_table_482_1_sva_dfm_1 = sigmoid_table_482_1_sva | (~ initialized_sva);
  assign sigmoid_table_536_1_sva_dfm_1 = sigmoid_table_536_1_sva | (~ initialized_sva);
  assign sigmoid_table_537_1_sva_dfm_1 = sigmoid_table_537_1_sva | (~ initialized_sva);
  assign sigmoid_table_538_1_sva_dfm_1 = sigmoid_table_538_1_sva | (~ initialized_sva);
  assign sigmoid_table_539_1_sva_dfm_1 = sigmoid_table_539_1_sva | (~ initialized_sva);
  assign sigmoid_table_540_1_sva_dfm_1 = sigmoid_table_540_1_sva | (~ initialized_sva);
  assign sigmoid_table_541_1_sva_dfm_1 = sigmoid_table_541_1_sva | (~ initialized_sva);
  assign sigmoid_table_552_1_sva_dfm_1 = sigmoid_table_552_1_sva | (~ initialized_sva);
  assign sigmoid_table_553_1_sva_dfm_1 = sigmoid_table_553_1_sva | (~ initialized_sva);
  assign sigmoid_table_554_1_sva_dfm_1 = sigmoid_table_554_1_sva | (~ initialized_sva);
  assign sigmoid_table_561_1_sva_dfm_1 = sigmoid_table_561_1_sva | (~ initialized_sva);
  assign sigmoid_table_562_1_sva_dfm_1 = sigmoid_table_562_1_sva | (~ initialized_sva);
  assign sigmoid_table_568_1_sva_dfm_1 = sigmoid_table_568_1_sva | (~ initialized_sva);
  assign sigmoid_table_569_1_sva_dfm_1 = sigmoid_table_569_1_sva | (~ initialized_sva);
  assign sigmoid_table_574_1_sva_dfm_1 = sigmoid_table_574_1_sva | (~ initialized_sva);
  assign sigmoid_table_578_1_sva_dfm_1 = sigmoid_table_578_1_sva | (~ initialized_sva);
  assign sigmoid_table_583_1_sva_dfm_1 = sigmoid_table_583_1_sva | (~ initialized_sva);
  assign sigmoid_table_586_1_sva_dfm_1 = sigmoid_table_586_1_sva | (~ initialized_sva);
  assign sigmoid_table_590_1_sva_dfm_1 = sigmoid_table_590_1_sva | (~ initialized_sva);
  assign sigmoid_table_593_1_sva_dfm_1 = sigmoid_table_593_1_sva | (~ initialized_sva);
  assign sigmoid_table_596_1_sva_dfm_1 = sigmoid_table_596_1_sva | (~ initialized_sva);
  assign sigmoid_table_599_1_sva_dfm_1 = sigmoid_table_599_1_sva | (~ initialized_sva);
  assign sigmoid_table_602_1_sva_dfm_1 = sigmoid_table_602_1_sva | (~ initialized_sva);
  assign sigmoid_table_607_1_sva_dfm_1 = sigmoid_table_607_1_sva | (~ initialized_sva);
  assign sigmoid_table_612_1_sva_dfm_1 = sigmoid_table_612_1_sva | (~ initialized_sva);
  assign sigmoid_table_619_1_sva_dfm_1 = sigmoid_table_619_1_sva | (~ initialized_sva);
  assign sigmoid_table_621_1_sva_dfm_1 = sigmoid_table_621_1_sva | (~ initialized_sva);
  assign sigmoid_table_623_1_sva_dfm_1 = sigmoid_table_623_1_sva | (~ initialized_sva);
  assign sigmoid_table_625_1_sva_dfm_1 = sigmoid_table_625_1_sva | (~ initialized_sva);
  assign sigmoid_table_627_1_sva_dfm_1 = sigmoid_table_627_1_sva | (~ initialized_sva);
  assign sigmoid_table_629_1_sva_dfm_1 = sigmoid_table_629_1_sva | (~ initialized_sva);
  assign sigmoid_table_638_1_sva_dfm_1 = sigmoid_table_638_1_sva | (~ initialized_sva);
  assign sigmoid_table_643_1_sva_dfm_1 = sigmoid_table_643_1_sva | (~ initialized_sva);
  assign sigmoid_table_645_1_sva_dfm_1 = sigmoid_table_645_1_sva | (~ initialized_sva);
  assign sigmoid_table_648_1_sva_dfm_1 = sigmoid_table_648_1_sva | (~ initialized_sva);
  assign sigmoid_table_653_1_sva_dfm_1 = sigmoid_table_653_1_sva | (~ initialized_sva);
  assign sigmoid_table_656_1_sva_dfm_1 = sigmoid_table_656_1_sva | (~ initialized_sva);
  assign sigmoid_table_659_1_sva_dfm_1 = sigmoid_table_659_1_sva | (~ initialized_sva);
  assign sigmoid_table_662_1_sva_dfm_1 = sigmoid_table_662_1_sva | (~ initialized_sva);
  assign sigmoid_table_665_1_sva_dfm_1 = sigmoid_table_665_1_sva | (~ initialized_sva);
  assign sigmoid_table_669_1_sva_dfm_1 = sigmoid_table_669_1_sva | (~ initialized_sva);
  assign sigmoid_table_672_1_sva_dfm_1 = sigmoid_table_672_1_sva | (~ initialized_sva);
  assign sigmoid_table_676_1_sva_dfm_1 = sigmoid_table_676_1_sva | (~ initialized_sva);
  assign sigmoid_table_680_1_sva_dfm_1 = sigmoid_table_680_1_sva | (~ initialized_sva);
  assign sigmoid_table_684_1_sva_dfm_1 = sigmoid_table_684_1_sva | (~ initialized_sva);
  assign sigmoid_table_688_1_sva_dfm_1 = sigmoid_table_688_1_sva | (~ initialized_sva);
  assign sigmoid_table_693_1_sva_dfm_1 = sigmoid_table_693_1_sva | (~ initialized_sva);
  assign sigmoid_table_697_1_sva_dfm_1 = sigmoid_table_697_1_sva | (~ initialized_sva);
  assign sigmoid_table_698_1_sva_dfm_1 = sigmoid_table_698_1_sva | (~ initialized_sva);
  assign sigmoid_table_703_1_sva_dfm_1 = sigmoid_table_703_1_sva | (~ initialized_sva);
  assign sigmoid_table_708_1_sva_dfm_1 = sigmoid_table_708_1_sva | (~ initialized_sva);
  assign sigmoid_table_709_1_sva_dfm_1 = sigmoid_table_709_1_sva | (~ initialized_sva);
  assign sigmoid_table_714_1_sva_dfm_1 = sigmoid_table_714_1_sva | (~ initialized_sva);
  assign sigmoid_table_715_1_sva_dfm_1 = sigmoid_table_715_1_sva | (~ initialized_sva);
  assign sigmoid_table_721_1_sva_dfm_1 = sigmoid_table_721_1_sva | (~ initialized_sva);
  assign sigmoid_table_722_1_sva_dfm_1 = sigmoid_table_722_1_sva | (~ initialized_sva);
  assign sigmoid_table_728_1_sva_dfm_1 = sigmoid_table_728_1_sva | (~ initialized_sva);
  assign sigmoid_table_729_1_sva_dfm_1 = sigmoid_table_729_1_sva | (~ initialized_sva);
  assign sigmoid_table_737_1_sva_dfm_1 = sigmoid_table_737_1_sva | (~ initialized_sva);
  assign sigmoid_table_738_1_sva_dfm_1 = sigmoid_table_738_1_sva | (~ initialized_sva);
  assign sigmoid_table_746_1_sva_dfm_1 = sigmoid_table_746_1_sva | (~ initialized_sva);
  assign sigmoid_table_747_1_sva_dfm_1 = sigmoid_table_747_1_sva | (~ initialized_sva);
  assign sigmoid_table_757_1_sva_dfm_1 = sigmoid_table_757_1_sva | (~ initialized_sva);
  assign sigmoid_table_758_1_sva_dfm_1 = sigmoid_table_758_1_sva | (~ initialized_sva);
  assign sigmoid_table_759_1_sva_dfm_1 = sigmoid_table_759_1_sva | (~ initialized_sva);
  assign sigmoid_table_770_1_sva_dfm_1 = sigmoid_table_770_1_sva | (~ initialized_sva);
  assign sigmoid_table_771_1_sva_dfm_1 = sigmoid_table_771_1_sva | (~ initialized_sva);
  assign sigmoid_table_772_1_sva_dfm_1 = sigmoid_table_772_1_sva | (~ initialized_sva);
  assign sigmoid_table_773_1_sva_dfm_1 = sigmoid_table_773_1_sva | (~ initialized_sva);
  assign sigmoid_table_786_1_sva_dfm_1 = sigmoid_table_786_1_sva | (~ initialized_sva);
  assign sigmoid_table_787_1_sva_dfm_1 = sigmoid_table_787_1_sva | (~ initialized_sva);
  assign sigmoid_table_788_1_sva_dfm_1 = sigmoid_table_788_1_sva | (~ initialized_sva);
  assign sigmoid_table_789_1_sva_dfm_1 = sigmoid_table_789_1_sva | (~ initialized_sva);
  assign sigmoid_table_790_1_sva_dfm_1 = sigmoid_table_790_1_sva | (~ initialized_sva);
  assign sigmoid_table_808_1_sva_dfm_1 = sigmoid_table_808_1_sva | (~ initialized_sva);
  assign sigmoid_table_809_1_sva_dfm_1 = sigmoid_table_809_1_sva | (~ initialized_sva);
  assign sigmoid_table_810_1_sva_dfm_1 = sigmoid_table_810_1_sva | (~ initialized_sva);
  assign sigmoid_table_811_1_sva_dfm_1 = sigmoid_table_811_1_sva | (~ initialized_sva);
  assign sigmoid_table_812_1_sva_dfm_1 = sigmoid_table_812_1_sva | (~ initialized_sva);
  assign sigmoid_table_813_1_sva_dfm_1 = sigmoid_table_813_1_sva | (~ initialized_sva);
  assign sigmoid_table_814_1_sva_dfm_1 = sigmoid_table_814_1_sva | (~ initialized_sva);
  assign sigmoid_table_841_1_sva_dfm_1 = sigmoid_table_841_1_sva | (~ initialized_sva);
  assign sigmoid_table_842_1_sva_dfm_1 = sigmoid_table_842_1_sva | (~ initialized_sva);
  assign sigmoid_table_843_1_sva_dfm_1 = sigmoid_table_843_1_sva | (~ initialized_sva);
  assign sigmoid_table_844_1_sva_dfm_1 = sigmoid_table_844_1_sva | (~ initialized_sva);
  assign sigmoid_table_845_1_sva_dfm_1 = sigmoid_table_845_1_sva | (~ initialized_sva);
  assign sigmoid_table_846_1_sva_dfm_1 = sigmoid_table_846_1_sva | (~ initialized_sva);
  assign sigmoid_table_847_1_sva_dfm_1 = sigmoid_table_847_1_sva | (~ initialized_sva);
  assign sigmoid_table_848_1_sva_dfm_1 = sigmoid_table_848_1_sva | (~ initialized_sva);
  assign sigmoid_table_849_1_sva_dfm_1 = sigmoid_table_849_1_sva | (~ initialized_sva);
  assign sigmoid_table_850_1_sva_dfm_1 = sigmoid_table_850_1_sva | (~ initialized_sva);
  assign sigmoid_table_851_1_sva_dfm_1 = sigmoid_table_851_1_sva | (~ initialized_sva);
  assign sigmoid_table_852_1_sva_dfm_1 = sigmoid_table_852_1_sva | (~ initialized_sva);
  assign sigmoid_table_442_8_sva_dfm_1 = sigmoid_table_442_8_sva | (~ initialized_sva);
  assign sigmoid_table_443_8_sva_dfm_1 = sigmoid_table_443_8_sva | (~ initialized_sva);
  assign sigmoid_table_444_8_sva_dfm_1 = sigmoid_table_444_8_sva | (~ initialized_sva);
  assign sigmoid_table_445_8_sva_dfm_1 = sigmoid_table_445_8_sva | (~ initialized_sva);
  assign sigmoid_table_446_8_sva_dfm_1 = sigmoid_table_446_8_sva | (~ initialized_sva);
  assign sigmoid_table_447_8_sva_dfm_1 = sigmoid_table_447_8_sva | (~ initialized_sva);
  assign sigmoid_table_448_8_sva_dfm_1 = sigmoid_table_448_8_sva | (~ initialized_sva);
  assign sigmoid_table_449_8_sva_dfm_1 = sigmoid_table_449_8_sva | (~ initialized_sva);
  assign sigmoid_table_450_8_sva_dfm_1 = sigmoid_table_450_8_sva | (~ initialized_sva);
  assign sigmoid_table_451_8_sva_dfm_1 = sigmoid_table_451_8_sva | (~ initialized_sva);
  assign sigmoid_table_452_8_sva_dfm_1 = sigmoid_table_452_8_sva | (~ initialized_sva);
  assign sigmoid_table_453_8_sva_dfm_1 = sigmoid_table_453_8_sva | (~ initialized_sva);
  assign sigmoid_table_454_8_sva_dfm_1 = sigmoid_table_454_8_sva | (~ initialized_sva);
  assign sigmoid_table_455_8_sva_dfm_1 = sigmoid_table_455_8_sva | (~ initialized_sva);
  assign sigmoid_table_456_8_sva_dfm_1 = sigmoid_table_456_8_sva | (~ initialized_sva);
  assign sigmoid_table_457_8_sva_dfm_1 = sigmoid_table_457_8_sva | (~ initialized_sva);
  assign sigmoid_table_458_8_sva_dfm_1 = sigmoid_table_458_8_sva | (~ initialized_sva);
  assign sigmoid_table_459_8_sva_dfm_1 = sigmoid_table_459_8_sva | (~ initialized_sva);
  assign sigmoid_table_460_8_sva_dfm_1 = sigmoid_table_460_8_sva | (~ initialized_sva);
  assign sigmoid_table_461_8_sva_dfm_1 = sigmoid_table_461_8_sva | (~ initialized_sva);
  assign sigmoid_table_462_8_sva_dfm_1 = sigmoid_table_462_8_sva | (~ initialized_sva);
  assign sigmoid_table_463_8_sva_dfm_1 = sigmoid_table_463_8_sva | (~ initialized_sva);
  assign sigmoid_table_464_8_sva_dfm_1 = sigmoid_table_464_8_sva | (~ initialized_sva);
  assign sigmoid_table_465_8_sva_dfm_1 = sigmoid_table_465_8_sva | (~ initialized_sva);
  assign sigmoid_table_466_8_sva_dfm_1 = sigmoid_table_466_8_sva | (~ initialized_sva);
  assign sigmoid_table_467_8_sva_dfm_1 = sigmoid_table_467_8_sva | (~ initialized_sva);
  assign sigmoid_table_468_8_sva_dfm_1 = sigmoid_table_468_8_sva | (~ initialized_sva);
  assign sigmoid_table_469_8_sva_dfm_1 = sigmoid_table_469_8_sva | (~ initialized_sva);
  assign sigmoid_table_470_8_sva_dfm_1 = sigmoid_table_470_8_sva | (~ initialized_sva);
  assign sigmoid_table_471_8_sva_dfm_1 = sigmoid_table_471_8_sva | (~ initialized_sva);
  assign sigmoid_table_472_8_sva_dfm_1 = sigmoid_table_472_8_sva | (~ initialized_sva);
  assign sigmoid_table_473_8_sva_dfm_1 = sigmoid_table_473_8_sva | (~ initialized_sva);
  assign sigmoid_table_474_8_sva_dfm_1 = sigmoid_table_474_8_sva | (~ initialized_sva);
  assign sigmoid_table_475_8_sva_dfm_1 = sigmoid_table_475_8_sva | (~ initialized_sva);
  assign sigmoid_table_476_8_sva_dfm_1 = sigmoid_table_476_8_sva | (~ initialized_sva);
  assign sigmoid_table_477_8_sva_dfm_1 = sigmoid_table_477_8_sva | (~ initialized_sva);
  assign sigmoid_table_478_8_sva_dfm_1 = sigmoid_table_478_8_sva | (~ initialized_sva);
  assign sigmoid_table_479_8_sva_dfm_1 = sigmoid_table_479_8_sva | (~ initialized_sva);
  assign sigmoid_table_480_7_sva_dfm_1 = sigmoid_table_480_7_sva | (~ initialized_sva);
  assign sigmoid_table_481_7_sva_dfm_1 = sigmoid_table_481_7_sva | (~ initialized_sva);
  assign sigmoid_table_482_7_sva_dfm_1 = sigmoid_table_482_7_sva | (~ initialized_sva);
  assign sigmoid_table_483_7_sva_dfm_1 = sigmoid_table_483_7_sva | (~ initialized_sva);
  assign sigmoid_table_484_7_sva_dfm_1 = sigmoid_table_484_7_sva | (~ initialized_sva);
  assign sigmoid_table_485_7_sva_dfm_1 = sigmoid_table_485_7_sva | (~ initialized_sva);
  assign sigmoid_table_486_7_sva_dfm_1 = sigmoid_table_486_7_sva | (~ initialized_sva);
  assign sigmoid_table_487_7_sva_dfm_1 = sigmoid_table_487_7_sva | (~ initialized_sva);
  assign sigmoid_table_488_7_sva_dfm_1 = sigmoid_table_488_7_sva | (~ initialized_sva);
  assign sigmoid_table_489_7_sva_dfm_1 = sigmoid_table_489_7_sva | (~ initialized_sva);
  assign sigmoid_table_490_7_sva_dfm_1 = sigmoid_table_490_7_sva | (~ initialized_sva);
  assign sigmoid_table_491_7_sva_dfm_1 = sigmoid_table_491_7_sva | (~ initialized_sva);
  assign sigmoid_table_492_7_sva_dfm_1 = sigmoid_table_492_7_sva | (~ initialized_sva);
  assign sigmoid_table_493_7_sva_dfm_1 = sigmoid_table_493_7_sva | (~ initialized_sva);
  assign sigmoid_table_494_7_sva_dfm_1 = sigmoid_table_494_7_sva | (~ initialized_sva);
  assign sigmoid_table_495_7_sva_dfm_1 = sigmoid_table_495_7_sva | (~ initialized_sva);
  assign sigmoid_table_496_6_sva_dfm_1 = sigmoid_table_496_6_sva | (~ initialized_sva);
  assign sigmoid_table_497_6_sva_dfm_1 = sigmoid_table_497_6_sva | (~ initialized_sva);
  assign sigmoid_table_498_6_sva_dfm_1 = sigmoid_table_498_6_sva | (~ initialized_sva);
  assign sigmoid_table_499_6_sva_dfm_1 = sigmoid_table_499_6_sva | (~ initialized_sva);
  assign sigmoid_table_500_6_sva_dfm_1 = sigmoid_table_500_6_sva | (~ initialized_sva);
  assign sigmoid_table_501_6_sva_dfm_1 = sigmoid_table_501_6_sva | (~ initialized_sva);
  assign sigmoid_table_502_6_sva_dfm_1 = sigmoid_table_502_6_sva | (~ initialized_sva);
  assign sigmoid_table_503_6_sva_dfm_1 = sigmoid_table_503_6_sva | (~ initialized_sva);
  assign sigmoid_table_504_5_sva_dfm_1 = sigmoid_table_504_5_sva | (~ initialized_sva);
  assign sigmoid_table_505_5_sva_dfm_1 = sigmoid_table_505_5_sva | (~ initialized_sva);
  assign sigmoid_table_506_5_sva_dfm_1 = sigmoid_table_506_5_sva | (~ initialized_sva);
  assign sigmoid_table_507_5_sva_dfm_1 = sigmoid_table_507_5_sva | (~ initialized_sva);
  assign sigmoid_table_508_4_sva_dfm_1 = sigmoid_table_508_4_sva | (~ initialized_sva);
  assign sigmoid_table_509_4_sva_dfm_1 = sigmoid_table_509_4_sva | (~ initialized_sva);
  assign sigmoid_table_510_3_sva_dfm_1 = sigmoid_table_510_3_sva | (~ initialized_sva);
  assign sigmoid_table_511_2_sva_dfm_1 = sigmoid_table_511_2_sva | (~ initialized_sva);
  assign sigmoid_table_158_2_sva_dfm_1 = sigmoid_table_158_2_sva | (~ initialized_sva);
  assign sigmoid_table_159_2_sva_dfm_1 = sigmoid_table_159_2_sva | (~ initialized_sva);
  assign sigmoid_table_160_2_sva_dfm_1 = sigmoid_table_160_2_sva | (~ initialized_sva);
  assign sigmoid_table_161_2_sva_dfm_1 = sigmoid_table_161_2_sva | (~ initialized_sva);
  assign sigmoid_table_162_2_sva_dfm_1 = sigmoid_table_162_2_sva | (~ initialized_sva);
  assign sigmoid_table_163_2_sva_dfm_1 = sigmoid_table_163_2_sva | (~ initialized_sva);
  assign sigmoid_table_164_2_sva_dfm_1 = sigmoid_table_164_2_sva | (~ initialized_sva);
  assign sigmoid_table_165_2_sva_dfm_1 = sigmoid_table_165_2_sva | (~ initialized_sva);
  assign sigmoid_table_166_2_sva_dfm_1 = sigmoid_table_166_2_sva | (~ initialized_sva);
  assign sigmoid_table_167_2_sva_dfm_1 = sigmoid_table_167_2_sva | (~ initialized_sva);
  assign sigmoid_table_168_2_sva_dfm_1 = sigmoid_table_168_2_sva | (~ initialized_sva);
  assign sigmoid_table_169_2_sva_dfm_1 = sigmoid_table_169_2_sva | (~ initialized_sva);
  assign sigmoid_table_170_2_sva_dfm_1 = sigmoid_table_170_2_sva | (~ initialized_sva);
  assign sigmoid_table_171_2_sva_dfm_1 = sigmoid_table_171_2_sva | (~ initialized_sva);
  assign sigmoid_table_172_2_sva_dfm_1 = sigmoid_table_172_2_sva | (~ initialized_sva);
  assign sigmoid_table_173_2_sva_dfm_1 = sigmoid_table_173_2_sva | (~ initialized_sva);
  assign sigmoid_table_174_2_sva_dfm_1 = sigmoid_table_174_2_sva | (~ initialized_sva);
  assign sigmoid_table_175_2_sva_dfm_1 = sigmoid_table_175_2_sva | (~ initialized_sva);
  assign sigmoid_table_176_2_sva_dfm_1 = sigmoid_table_176_2_sva | (~ initialized_sva);
  assign sigmoid_table_177_2_sva_dfm_1 = sigmoid_table_177_2_sva | (~ initialized_sva);
  assign sigmoid_table_178_2_sva_dfm_1 = sigmoid_table_178_2_sva | (~ initialized_sva);
  assign sigmoid_table_179_2_sva_dfm_1 = sigmoid_table_179_2_sva | (~ initialized_sva);
  assign sigmoid_table_180_2_sva_dfm_1 = sigmoid_table_180_2_sva | (~ initialized_sva);
  assign sigmoid_table_181_2_sva_dfm_1 = sigmoid_table_181_2_sva | (~ initialized_sva);
  assign sigmoid_table_182_2_sva_dfm_1 = sigmoid_table_182_2_sva | (~ initialized_sva);
  assign sigmoid_table_183_2_sva_dfm_1 = sigmoid_table_183_2_sva | (~ initialized_sva);
  assign sigmoid_table_229_2_sva_dfm_1 = sigmoid_table_229_2_sva | (~ initialized_sva);
  assign sigmoid_table_230_2_sva_dfm_1 = sigmoid_table_230_2_sva | (~ initialized_sva);
  assign sigmoid_table_231_2_sva_dfm_1 = sigmoid_table_231_2_sva | (~ initialized_sva);
  assign sigmoid_table_232_2_sva_dfm_1 = sigmoid_table_232_2_sva | (~ initialized_sva);
  assign sigmoid_table_233_2_sva_dfm_1 = sigmoid_table_233_2_sva | (~ initialized_sva);
  assign sigmoid_table_234_2_sva_dfm_1 = sigmoid_table_234_2_sva | (~ initialized_sva);
  assign sigmoid_table_235_2_sva_dfm_1 = sigmoid_table_235_2_sva | (~ initialized_sva);
  assign sigmoid_table_236_2_sva_dfm_1 = sigmoid_table_236_2_sva | (~ initialized_sva);
  assign sigmoid_table_237_2_sva_dfm_1 = sigmoid_table_237_2_sva | (~ initialized_sva);
  assign sigmoid_table_238_2_sva_dfm_1 = sigmoid_table_238_2_sva | (~ initialized_sva);
  assign sigmoid_table_262_2_sva_dfm_1 = sigmoid_table_262_2_sva | (~ initialized_sva);
  assign sigmoid_table_263_2_sva_dfm_1 = sigmoid_table_263_2_sva | (~ initialized_sva);
  assign sigmoid_table_264_2_sva_dfm_1 = sigmoid_table_264_2_sva | (~ initialized_sva);
  assign sigmoid_table_265_2_sva_dfm_1 = sigmoid_table_265_2_sva | (~ initialized_sva);
  assign sigmoid_table_266_2_sva_dfm_1 = sigmoid_table_266_2_sva | (~ initialized_sva);
  assign sigmoid_table_267_2_sva_dfm_1 = sigmoid_table_267_2_sva | (~ initialized_sva);
  assign sigmoid_table_284_2_sva_dfm_1 = sigmoid_table_284_2_sva | (~ initialized_sva);
  assign sigmoid_table_285_2_sva_dfm_1 = sigmoid_table_285_2_sva | (~ initialized_sva);
  assign sigmoid_table_286_2_sva_dfm_1 = sigmoid_table_286_2_sva | (~ initialized_sva);
  assign sigmoid_table_287_2_sva_dfm_1 = sigmoid_table_287_2_sva | (~ initialized_sva);
  assign sigmoid_table_301_2_sva_dfm_1 = sigmoid_table_301_2_sva | (~ initialized_sva);
  assign sigmoid_table_302_2_sva_dfm_1 = sigmoid_table_302_2_sva | (~ initialized_sva);
  assign sigmoid_table_303_2_sva_dfm_1 = sigmoid_table_303_2_sva | (~ initialized_sva);
  assign sigmoid_table_314_2_sva_dfm_1 = sigmoid_table_314_2_sva | (~ initialized_sva);
  assign sigmoid_table_315_2_sva_dfm_1 = sigmoid_table_315_2_sva | (~ initialized_sva);
  assign sigmoid_table_316_2_sva_dfm_1 = sigmoid_table_316_2_sva | (~ initialized_sva);
  assign sigmoid_table_325_2_sva_dfm_1 = sigmoid_table_325_2_sva | (~ initialized_sva);
  assign sigmoid_table_326_2_sva_dfm_1 = sigmoid_table_326_2_sva | (~ initialized_sva);
  assign sigmoid_table_327_2_sva_dfm_1 = sigmoid_table_327_2_sva | (~ initialized_sva);
  assign sigmoid_table_335_2_sva_dfm_1 = sigmoid_table_335_2_sva | (~ initialized_sva);
  assign sigmoid_table_336_2_sva_dfm_1 = sigmoid_table_336_2_sva | (~ initialized_sva);
  assign sigmoid_table_343_2_sva_dfm_1 = sigmoid_table_343_2_sva | (~ initialized_sva);
  assign sigmoid_table_344_2_sva_dfm_1 = sigmoid_table_344_2_sva | (~ initialized_sva);
  assign sigmoid_table_351_2_sva_dfm_1 = sigmoid_table_351_2_sva | (~ initialized_sva);
  assign sigmoid_table_352_2_sva_dfm_1 = sigmoid_table_352_2_sva | (~ initialized_sva);
  assign sigmoid_table_358_2_sva_dfm_1 = sigmoid_table_358_2_sva | (~ initialized_sva);
  assign sigmoid_table_359_2_sva_dfm_1 = sigmoid_table_359_2_sva | (~ initialized_sva);
  assign sigmoid_table_364_2_sva_dfm_1 = sigmoid_table_364_2_sva | (~ initialized_sva);
  assign sigmoid_table_365_2_sva_dfm_1 = sigmoid_table_365_2_sva | (~ initialized_sva);
  assign sigmoid_table_370_2_sva_dfm_1 = sigmoid_table_370_2_sva | (~ initialized_sva);
  assign sigmoid_table_371_2_sva_dfm_1 = sigmoid_table_371_2_sva | (~ initialized_sva);
  assign sigmoid_table_376_2_sva_dfm_1 = sigmoid_table_376_2_sva | (~ initialized_sva);
  assign sigmoid_table_381_2_sva_dfm_1 = sigmoid_table_381_2_sva | (~ initialized_sva);
  assign sigmoid_table_386_2_sva_dfm_1 = sigmoid_table_386_2_sva | (~ initialized_sva);
  assign sigmoid_table_390_2_sva_dfm_1 = sigmoid_table_390_2_sva | (~ initialized_sva);
  assign sigmoid_table_395_2_sva_dfm_1 = sigmoid_table_395_2_sva | (~ initialized_sva);
  assign sigmoid_table_399_2_sva_dfm_1 = sigmoid_table_399_2_sva | (~ initialized_sva);
  assign sigmoid_table_403_2_sva_dfm_1 = sigmoid_table_403_2_sva | (~ initialized_sva);
  assign sigmoid_table_406_2_sva_dfm_1 = sigmoid_table_406_2_sva | (~ initialized_sva);
  assign sigmoid_table_410_2_sva_dfm_1 = sigmoid_table_410_2_sva | (~ initialized_sva);
  assign sigmoid_table_417_2_sva_dfm_1 = sigmoid_table_417_2_sva | (~ initialized_sva);
  assign sigmoid_table_420_2_sva_dfm_1 = sigmoid_table_420_2_sva | (~ initialized_sva);
  assign sigmoid_table_423_2_sva_dfm_1 = sigmoid_table_423_2_sva | (~ initialized_sva);
  assign sigmoid_table_432_2_sva_dfm_1 = sigmoid_table_432_2_sva | (~ initialized_sva);
  assign sigmoid_table_435_2_sva_dfm_1 = sigmoid_table_435_2_sva | (~ initialized_sva);
  assign sigmoid_table_438_2_sva_dfm_1 = sigmoid_table_438_2_sva | (~ initialized_sva);
  assign sigmoid_table_441_2_sva_dfm_1 = sigmoid_table_441_2_sva | (~ initialized_sva);
  assign sigmoid_table_446_2_sva_dfm_1 = sigmoid_table_446_2_sva | (~ initialized_sva);
  assign sigmoid_table_451_2_sva_dfm_1 = sigmoid_table_451_2_sva | (~ initialized_sva);
  assign sigmoid_table_456_2_sva_dfm_1 = sigmoid_table_456_2_sva | (~ initialized_sva);
  assign sigmoid_table_463_2_sva_dfm_1 = sigmoid_table_463_2_sva | (~ initialized_sva);
  assign sigmoid_table_465_2_sva_dfm_1 = sigmoid_table_465_2_sva | (~ initialized_sva);
  assign sigmoid_table_470_2_sva_dfm_1 = sigmoid_table_470_2_sva | (~ initialized_sva);
  assign sigmoid_table_472_2_sva_dfm_1 = sigmoid_table_472_2_sva | (~ initialized_sva);
  assign sigmoid_table_474_2_sva_dfm_1 = sigmoid_table_474_2_sva | (~ initialized_sva);
  assign sigmoid_table_483_2_sva_dfm_1 = sigmoid_table_483_2_sva | (~ initialized_sva);
  assign sigmoid_table_485_2_sva_dfm_1 = sigmoid_table_485_2_sva | (~ initialized_sva);
  assign sigmoid_table_487_2_sva_dfm_1 = sigmoid_table_487_2_sva | (~ initialized_sva);
  assign sigmoid_table_489_2_sva_dfm_1 = sigmoid_table_489_2_sva | (~ initialized_sva);
  assign sigmoid_table_491_2_sva_dfm_1 = sigmoid_table_491_2_sva | (~ initialized_sva);
  assign sigmoid_table_493_2_sva_dfm_1 = sigmoid_table_493_2_sva | (~ initialized_sva);
  assign sigmoid_table_495_2_sva_dfm_1 = sigmoid_table_495_2_sva | (~ initialized_sva);
  assign sigmoid_table_497_2_sva_dfm_1 = sigmoid_table_497_2_sva | (~ initialized_sva);
  assign sigmoid_table_499_2_sva_dfm_1 = sigmoid_table_499_2_sva | (~ initialized_sva);
  assign sigmoid_table_501_2_sva_dfm_1 = sigmoid_table_501_2_sva | (~ initialized_sva);
  assign sigmoid_table_503_2_sva_dfm_1 = sigmoid_table_503_2_sva | (~ initialized_sva);
  assign sigmoid_table_505_2_sva_dfm_1 = sigmoid_table_505_2_sva | (~ initialized_sva);
  assign sigmoid_table_507_2_sva_dfm_1 = sigmoid_table_507_2_sva | (~ initialized_sva);
  assign sigmoid_table_509_2_sva_dfm_1 = sigmoid_table_509_2_sva | (~ initialized_sva);
  assign sigmoid_table_513_2_sva_dfm_1 = sigmoid_table_513_2_sva | (~ initialized_sva);
  assign sigmoid_table_515_2_sva_dfm_1 = sigmoid_table_515_2_sva | (~ initialized_sva);
  assign sigmoid_table_542_2_sva_dfm_1 = sigmoid_table_542_2_sva | (~ initialized_sva);
  assign sigmoid_table_544_2_sva_dfm_1 = sigmoid_table_544_2_sva | (~ initialized_sva);
  assign sigmoid_table_546_2_sva_dfm_1 = sigmoid_table_546_2_sva | (~ initialized_sva);
  assign sigmoid_table_548_2_sva_dfm_1 = sigmoid_table_548_2_sva | (~ initialized_sva);
  assign sigmoid_table_555_2_sva_dfm_1 = sigmoid_table_555_2_sva | (~ initialized_sva);
  assign sigmoid_table_557_2_sva_dfm_1 = sigmoid_table_557_2_sva | (~ initialized_sva);
  assign sigmoid_table_564_2_sva_dfm_1 = sigmoid_table_564_2_sva | (~ initialized_sva);
  assign sigmoid_table_566_2_sva_dfm_1 = sigmoid_table_566_2_sva | (~ initialized_sva);
  assign sigmoid_table_571_2_sva_dfm_1 = sigmoid_table_571_2_sva | (~ initialized_sva);
  assign sigmoid_table_576_2_sva_dfm_1 = sigmoid_table_576_2_sva | (~ initialized_sva);
  assign sigmoid_table_579_2_sva_dfm_1 = sigmoid_table_579_2_sva | (~ initialized_sva);
  assign sigmoid_table_581_2_sva_dfm_1 = sigmoid_table_581_2_sva | (~ initialized_sva);
  assign sigmoid_table_584_2_sva_dfm_1 = sigmoid_table_584_2_sva | (~ initialized_sva);
  assign sigmoid_table_587_2_sva_dfm_1 = sigmoid_table_587_2_sva | (~ initialized_sva);
  assign sigmoid_table_595_2_sva_dfm_1 = sigmoid_table_595_2_sva | (~ initialized_sva);
  assign sigmoid_table_598_2_sva_dfm_1 = sigmoid_table_598_2_sva | (~ initialized_sva);
  assign sigmoid_table_605_2_sva_dfm_1 = sigmoid_table_605_2_sva | (~ initialized_sva);
  assign sigmoid_table_608_2_sva_dfm_1 = sigmoid_table_608_2_sva | (~ initialized_sva);
  assign sigmoid_table_611_2_sva_dfm_1 = sigmoid_table_611_2_sva | (~ initialized_sva);
  assign sigmoid_table_615_2_sva_dfm_1 = sigmoid_table_615_2_sva | (~ initialized_sva);
  assign sigmoid_table_622_2_sva_dfm_1 = sigmoid_table_622_2_sva | (~ initialized_sva);
  assign sigmoid_table_626_2_sva_dfm_1 = sigmoid_table_626_2_sva | (~ initialized_sva);
  assign sigmoid_table_630_2_sva_dfm_1 = sigmoid_table_630_2_sva | (~ initialized_sva);
  assign sigmoid_table_631_2_sva_dfm_1 = sigmoid_table_631_2_sva | (~ initialized_sva);
  assign sigmoid_table_635_2_sva_dfm_1 = sigmoid_table_635_2_sva | (~ initialized_sva);
  assign sigmoid_table_639_2_sva_dfm_1 = sigmoid_table_639_2_sva | (~ initialized_sva);
  assign sigmoid_table_640_2_sva_dfm_1 = sigmoid_table_640_2_sva | (~ initialized_sva);
  assign sigmoid_table_644_2_sva_dfm_1 = sigmoid_table_644_2_sva | (~ initialized_sva);
  assign sigmoid_table_649_2_sva_dfm_1 = sigmoid_table_649_2_sva | (~ initialized_sva);
  assign sigmoid_table_650_2_sva_dfm_1 = sigmoid_table_650_2_sva | (~ initialized_sva);
  assign sigmoid_table_655_2_sva_dfm_1 = sigmoid_table_655_2_sva | (~ initialized_sva);
  assign sigmoid_table_661_2_sva_dfm_1 = sigmoid_table_661_2_sva | (~ initialized_sva);
  assign sigmoid_table_667_2_sva_dfm_1 = sigmoid_table_667_2_sva | (~ initialized_sva);
  assign sigmoid_table_668_2_sva_dfm_1 = sigmoid_table_668_2_sva | (~ initialized_sva);
  assign sigmoid_table_674_2_sva_dfm_1 = sigmoid_table_674_2_sva | (~ initialized_sva);
  assign sigmoid_table_675_2_sva_dfm_1 = sigmoid_table_675_2_sva | (~ initialized_sva);
  assign sigmoid_table_682_2_sva_dfm_1 = sigmoid_table_682_2_sva | (~ initialized_sva);
  assign sigmoid_table_683_2_sva_dfm_1 = sigmoid_table_683_2_sva | (~ initialized_sva);
  assign sigmoid_table_690_2_sva_dfm_1 = sigmoid_table_690_2_sva | (~ initialized_sva);
  assign sigmoid_table_691_2_sva_dfm_1 = sigmoid_table_691_2_sva | (~ initialized_sva);
  assign sigmoid_table_692_2_sva_dfm_1 = sigmoid_table_692_2_sva | (~ initialized_sva);
  assign sigmoid_table_700_2_sva_dfm_1 = sigmoid_table_700_2_sva | (~ initialized_sva);
  assign sigmoid_table_701_2_sva_dfm_1 = sigmoid_table_701_2_sva | (~ initialized_sva);
  assign sigmoid_table_702_2_sva_dfm_1 = sigmoid_table_702_2_sva | (~ initialized_sva);
  assign sigmoid_table_711_2_sva_dfm_1 = sigmoid_table_711_2_sva | (~ initialized_sva);
  assign sigmoid_table_712_2_sva_dfm_1 = sigmoid_table_712_2_sva | (~ initialized_sva);
  assign sigmoid_table_713_2_sva_dfm_1 = sigmoid_table_713_2_sva | (~ initialized_sva);
  assign sigmoid_table_724_2_sva_dfm_1 = sigmoid_table_724_2_sva | (~ initialized_sva);
  assign sigmoid_table_725_2_sva_dfm_1 = sigmoid_table_725_2_sva | (~ initialized_sva);
  assign sigmoid_table_726_2_sva_dfm_1 = sigmoid_table_726_2_sva | (~ initialized_sva);
  assign sigmoid_table_727_2_sva_dfm_1 = sigmoid_table_727_2_sva | (~ initialized_sva);
  assign sigmoid_table_741_2_sva_dfm_1 = sigmoid_table_741_2_sva | (~ initialized_sva);
  assign sigmoid_table_742_2_sva_dfm_1 = sigmoid_table_742_2_sva | (~ initialized_sva);
  assign sigmoid_table_743_2_sva_dfm_1 = sigmoid_table_743_2_sva | (~ initialized_sva);
  assign sigmoid_table_744_2_sva_dfm_1 = sigmoid_table_744_2_sva | (~ initialized_sva);
  assign sigmoid_table_745_2_sva_dfm_1 = sigmoid_table_745_2_sva | (~ initialized_sva);
  assign sigmoid_table_763_2_sva_dfm_1 = sigmoid_table_763_2_sva | (~ initialized_sva);
  assign sigmoid_table_764_2_sva_dfm_1 = sigmoid_table_764_2_sva | (~ initialized_sva);
  assign sigmoid_table_765_2_sva_dfm_1 = sigmoid_table_765_2_sva | (~ initialized_sva);
  assign sigmoid_table_766_2_sva_dfm_1 = sigmoid_table_766_2_sva | (~ initialized_sva);
  assign sigmoid_table_767_2_sva_dfm_1 = sigmoid_table_767_2_sva | (~ initialized_sva);
  assign sigmoid_table_768_2_sva_dfm_1 = sigmoid_table_768_2_sva | (~ initialized_sva);
  assign sigmoid_table_769_2_sva_dfm_1 = sigmoid_table_769_2_sva | (~ initialized_sva);
  assign sigmoid_table_796_2_sva_dfm_1 = sigmoid_table_796_2_sva | (~ initialized_sva);
  assign sigmoid_table_797_2_sva_dfm_1 = sigmoid_table_797_2_sva | (~ initialized_sva);
  assign sigmoid_table_798_2_sva_dfm_1 = sigmoid_table_798_2_sva | (~ initialized_sva);
  assign sigmoid_table_799_2_sva_dfm_1 = sigmoid_table_799_2_sva | (~ initialized_sva);
  assign sigmoid_table_800_2_sva_dfm_1 = sigmoid_table_800_2_sva | (~ initialized_sva);
  assign sigmoid_table_801_2_sva_dfm_1 = sigmoid_table_801_2_sva | (~ initialized_sva);
  assign sigmoid_table_802_2_sva_dfm_1 = sigmoid_table_802_2_sva | (~ initialized_sva);
  assign sigmoid_table_803_2_sva_dfm_1 = sigmoid_table_803_2_sva | (~ initialized_sva);
  assign sigmoid_table_804_2_sva_dfm_1 = sigmoid_table_804_2_sva | (~ initialized_sva);
  assign sigmoid_table_805_2_sva_dfm_1 = sigmoid_table_805_2_sva | (~ initialized_sva);
  assign sigmoid_table_806_2_sva_dfm_1 = sigmoid_table_806_2_sva | (~ initialized_sva);
  assign sigmoid_table_807_2_sva_dfm_1 = sigmoid_table_807_2_sva | (~ initialized_sva);
  assign sigmoid_table_388_7_sva_dfm_1 = sigmoid_table_388_7_sva | (~ initialized_sva);
  assign sigmoid_table_389_7_sva_dfm_1 = sigmoid_table_389_7_sva | (~ initialized_sva);
  assign sigmoid_table_390_7_sva_dfm_1 = sigmoid_table_390_7_sva | (~ initialized_sva);
  assign sigmoid_table_391_7_sva_dfm_1 = sigmoid_table_391_7_sva | (~ initialized_sva);
  assign sigmoid_table_392_7_sva_dfm_1 = sigmoid_table_392_7_sva | (~ initialized_sva);
  assign sigmoid_table_393_7_sva_dfm_1 = sigmoid_table_393_7_sva | (~ initialized_sva);
  assign sigmoid_table_394_7_sva_dfm_1 = sigmoid_table_394_7_sva | (~ initialized_sva);
  assign sigmoid_table_395_7_sva_dfm_1 = sigmoid_table_395_7_sva | (~ initialized_sva);
  assign sigmoid_table_396_7_sva_dfm_1 = sigmoid_table_396_7_sva | (~ initialized_sva);
  assign sigmoid_table_397_7_sva_dfm_1 = sigmoid_table_397_7_sva | (~ initialized_sva);
  assign sigmoid_table_398_7_sva_dfm_1 = sigmoid_table_398_7_sva | (~ initialized_sva);
  assign sigmoid_table_399_7_sva_dfm_1 = sigmoid_table_399_7_sva | (~ initialized_sva);
  assign sigmoid_table_400_7_sva_dfm_1 = sigmoid_table_400_7_sva | (~ initialized_sva);
  assign sigmoid_table_401_7_sva_dfm_1 = sigmoid_table_401_7_sva | (~ initialized_sva);
  assign sigmoid_table_402_7_sva_dfm_1 = sigmoid_table_402_7_sva | (~ initialized_sva);
  assign sigmoid_table_403_7_sva_dfm_1 = sigmoid_table_403_7_sva | (~ initialized_sva);
  assign sigmoid_table_404_7_sva_dfm_1 = sigmoid_table_404_7_sva | (~ initialized_sva);
  assign sigmoid_table_405_7_sva_dfm_1 = sigmoid_table_405_7_sva | (~ initialized_sva);
  assign sigmoid_table_406_7_sva_dfm_1 = sigmoid_table_406_7_sva | (~ initialized_sva);
  assign sigmoid_table_407_7_sva_dfm_1 = sigmoid_table_407_7_sva | (~ initialized_sva);
  assign sigmoid_table_408_7_sva_dfm_1 = sigmoid_table_408_7_sva | (~ initialized_sva);
  assign sigmoid_table_409_7_sva_dfm_1 = sigmoid_table_409_7_sva | (~ initialized_sva);
  assign sigmoid_table_410_7_sva_dfm_1 = sigmoid_table_410_7_sva | (~ initialized_sva);
  assign sigmoid_table_411_7_sva_dfm_1 = sigmoid_table_411_7_sva | (~ initialized_sva);
  assign sigmoid_table_412_7_sva_dfm_1 = sigmoid_table_412_7_sva | (~ initialized_sva);
  assign sigmoid_table_413_7_sva_dfm_1 = sigmoid_table_413_7_sva | (~ initialized_sva);
  assign sigmoid_table_414_7_sva_dfm_1 = sigmoid_table_414_7_sva | (~ initialized_sva);
  assign sigmoid_table_415_7_sva_dfm_1 = sigmoid_table_415_7_sva | (~ initialized_sva);
  assign sigmoid_table_416_7_sva_dfm_1 = sigmoid_table_416_7_sva | (~ initialized_sva);
  assign sigmoid_table_417_7_sva_dfm_1 = sigmoid_table_417_7_sva | (~ initialized_sva);
  assign sigmoid_table_418_7_sva_dfm_1 = sigmoid_table_418_7_sva | (~ initialized_sva);
  assign sigmoid_table_419_6_sva_dfm_1 = sigmoid_table_419_6_sva | (~ initialized_sva);
  assign sigmoid_table_420_6_sva_dfm_1 = sigmoid_table_420_6_sva | (~ initialized_sva);
  assign sigmoid_table_421_6_sva_dfm_1 = sigmoid_table_421_6_sva | (~ initialized_sva);
  assign sigmoid_table_422_6_sva_dfm_1 = sigmoid_table_422_6_sva | (~ initialized_sva);
  assign sigmoid_table_423_6_sva_dfm_1 = sigmoid_table_423_6_sva | (~ initialized_sva);
  assign sigmoid_table_424_6_sva_dfm_1 = sigmoid_table_424_6_sva | (~ initialized_sva);
  assign sigmoid_table_425_6_sva_dfm_1 = sigmoid_table_425_6_sva | (~ initialized_sva);
  assign sigmoid_table_426_6_sva_dfm_1 = sigmoid_table_426_6_sva | (~ initialized_sva);
  assign sigmoid_table_427_6_sva_dfm_1 = sigmoid_table_427_6_sva | (~ initialized_sva);
  assign sigmoid_table_428_6_sva_dfm_1 = sigmoid_table_428_6_sva | (~ initialized_sva);
  assign sigmoid_table_429_6_sva_dfm_1 = sigmoid_table_429_6_sva | (~ initialized_sva);
  assign sigmoid_table_430_6_sva_dfm_1 = sigmoid_table_430_6_sva | (~ initialized_sva);
  assign sigmoid_table_431_5_sva_dfm_1 = sigmoid_table_431_5_sva | (~ initialized_sva);
  assign sigmoid_table_432_5_sva_dfm_1 = sigmoid_table_432_5_sva | (~ initialized_sva);
  assign sigmoid_table_433_5_sva_dfm_1 = sigmoid_table_433_5_sva | (~ initialized_sva);
  assign sigmoid_table_434_5_sva_dfm_1 = sigmoid_table_434_5_sva | (~ initialized_sva);
  assign sigmoid_table_435_5_sva_dfm_1 = sigmoid_table_435_5_sva | (~ initialized_sva);
  assign sigmoid_table_436_5_sva_dfm_1 = sigmoid_table_436_5_sva | (~ initialized_sva);
  assign sigmoid_table_437_4_sva_dfm_1 = sigmoid_table_437_4_sva | (~ initialized_sva);
  assign sigmoid_table_438_4_sva_dfm_1 = sigmoid_table_438_4_sva | (~ initialized_sva);
  assign sigmoid_table_439_3_sva_dfm_1 = sigmoid_table_439_3_sva | (~ initialized_sva);
  assign sigmoid_table_440_3_sva_dfm_1 = sigmoid_table_440_3_sva | (~ initialized_sva);
  assign sigmoid_table_545_7_sva_dfm_1 = sigmoid_table_545_7_sva | (~ initialized_sva);
  assign sigmoid_table_546_7_sva_dfm_1 = sigmoid_table_546_7_sva | (~ initialized_sva);
  assign sigmoid_table_547_7_sva_dfm_1 = sigmoid_table_547_7_sva | (~ initialized_sva);
  assign sigmoid_table_548_7_sva_dfm_1 = sigmoid_table_548_7_sva | (~ initialized_sva);
  assign sigmoid_table_549_7_sva_dfm_1 = sigmoid_table_549_7_sva | (~ initialized_sva);
  assign sigmoid_table_550_7_sva_dfm_1 = sigmoid_table_550_7_sva | (~ initialized_sva);
  assign sigmoid_table_551_7_sva_dfm_1 = sigmoid_table_551_7_sva | (~ initialized_sva);
  assign sigmoid_table_552_7_sva_dfm_1 = sigmoid_table_552_7_sva | (~ initialized_sva);
  assign sigmoid_table_553_7_sva_dfm_1 = sigmoid_table_553_7_sva | (~ initialized_sva);
  assign sigmoid_table_554_7_sva_dfm_1 = sigmoid_table_554_7_sva | (~ initialized_sva);
  assign sigmoid_table_555_7_sva_dfm_1 = sigmoid_table_555_7_sva | (~ initialized_sva);
  assign sigmoid_table_556_7_sva_dfm_1 = sigmoid_table_556_7_sva | (~ initialized_sva);
  assign sigmoid_table_557_7_sva_dfm_1 = sigmoid_table_557_7_sva | (~ initialized_sva);
  assign sigmoid_table_558_7_sva_dfm_1 = sigmoid_table_558_7_sva | (~ initialized_sva);
  assign sigmoid_table_559_7_sva_dfm_1 = sigmoid_table_559_7_sva | (~ initialized_sva);
  assign sigmoid_table_560_7_sva_dfm_1 = sigmoid_table_560_7_sva | (~ initialized_sva);
  assign sigmoid_table_561_7_sva_dfm_1 = sigmoid_table_561_7_sva | (~ initialized_sva);
  assign sigmoid_table_562_7_sva_dfm_1 = sigmoid_table_562_7_sva | (~ initialized_sva);
  assign sigmoid_table_563_6_sva_dfm_1 = sigmoid_table_563_6_sva | (~ initialized_sva);
  assign sigmoid_table_564_6_sva_dfm_1 = sigmoid_table_564_6_sva | (~ initialized_sva);
  assign sigmoid_table_565_6_sva_dfm_1 = sigmoid_table_565_6_sva | (~ initialized_sva);
  assign sigmoid_table_566_6_sva_dfm_1 = sigmoid_table_566_6_sva | (~ initialized_sva);
  assign sigmoid_table_567_6_sva_dfm_1 = sigmoid_table_567_6_sva | (~ initialized_sva);
  assign sigmoid_table_568_6_sva_dfm_1 = sigmoid_table_568_6_sva | (~ initialized_sva);
  assign sigmoid_table_569_6_sva_dfm_1 = sigmoid_table_569_6_sva | (~ initialized_sva);
  assign sigmoid_table_570_6_sva_dfm_1 = sigmoid_table_570_6_sva | (~ initialized_sva);
  assign sigmoid_table_571_6_sva_dfm_1 = sigmoid_table_571_6_sva | (~ initialized_sva);
  assign sigmoid_table_572_6_sva_dfm_1 = sigmoid_table_572_6_sva | (~ initialized_sva);
  assign sigmoid_table_573_5_sva_dfm_1 = sigmoid_table_573_5_sva | (~ initialized_sva);
  assign sigmoid_table_574_5_sva_dfm_1 = sigmoid_table_574_5_sva | (~ initialized_sva);
  assign sigmoid_table_575_5_sva_dfm_1 = sigmoid_table_575_5_sva | (~ initialized_sva);
  assign sigmoid_table_576_5_sva_dfm_1 = sigmoid_table_576_5_sva | (~ initialized_sva);
  assign sigmoid_table_577_5_sva_dfm_1 = sigmoid_table_577_5_sva | (~ initialized_sva);
  assign sigmoid_table_578_4_sva_dfm_1 = sigmoid_table_578_4_sva | (~ initialized_sva);
  assign sigmoid_table_579_4_sva_dfm_1 = sigmoid_table_579_4_sva | (~ initialized_sva);
  assign sigmoid_table_580_3_sva_dfm_1 = sigmoid_table_580_3_sva | (~ initialized_sva);
  assign sigmoid_table_202_3_sva_dfm_1 = sigmoid_table_202_3_sva | (~ initialized_sva);
  assign sigmoid_table_203_3_sva_dfm_1 = sigmoid_table_203_3_sva | (~ initialized_sva);
  assign sigmoid_table_204_3_sva_dfm_1 = sigmoid_table_204_3_sva | (~ initialized_sva);
  assign sigmoid_table_205_3_sva_dfm_1 = sigmoid_table_205_3_sva | (~ initialized_sva);
  assign sigmoid_table_206_3_sva_dfm_1 = sigmoid_table_206_3_sva | (~ initialized_sva);
  assign sigmoid_table_207_3_sva_dfm_1 = sigmoid_table_207_3_sva | (~ initialized_sva);
  assign sigmoid_table_208_3_sva_dfm_1 = sigmoid_table_208_3_sva | (~ initialized_sva);
  assign sigmoid_table_209_3_sva_dfm_1 = sigmoid_table_209_3_sva | (~ initialized_sva);
  assign sigmoid_table_210_3_sva_dfm_1 = sigmoid_table_210_3_sva | (~ initialized_sva);
  assign sigmoid_table_211_3_sva_dfm_1 = sigmoid_table_211_3_sva | (~ initialized_sva);
  assign sigmoid_table_212_3_sva_dfm_1 = sigmoid_table_212_3_sva | (~ initialized_sva);
  assign sigmoid_table_213_3_sva_dfm_1 = sigmoid_table_213_3_sva | (~ initialized_sva);
  assign sigmoid_table_214_3_sva_dfm_1 = sigmoid_table_214_3_sva | (~ initialized_sva);
  assign sigmoid_table_215_3_sva_dfm_1 = sigmoid_table_215_3_sva | (~ initialized_sva);
  assign sigmoid_table_216_3_sva_dfm_1 = sigmoid_table_216_3_sva | (~ initialized_sva);
  assign sigmoid_table_217_3_sva_dfm_1 = sigmoid_table_217_3_sva | (~ initialized_sva);
  assign sigmoid_table_218_3_sva_dfm_1 = sigmoid_table_218_3_sva | (~ initialized_sva);
  assign sigmoid_table_219_3_sva_dfm_1 = sigmoid_table_219_3_sva | (~ initialized_sva);
  assign sigmoid_table_220_3_sva_dfm_1 = sigmoid_table_220_3_sva | (~ initialized_sva);
  assign sigmoid_table_221_3_sva_dfm_1 = sigmoid_table_221_3_sva | (~ initialized_sva);
  assign sigmoid_table_222_3_sva_dfm_1 = sigmoid_table_222_3_sva | (~ initialized_sva);
  assign sigmoid_table_223_3_sva_dfm_1 = sigmoid_table_223_3_sva | (~ initialized_sva);
  assign sigmoid_table_224_3_sva_dfm_1 = sigmoid_table_224_3_sva | (~ initialized_sva);
  assign sigmoid_table_225_3_sva_dfm_1 = sigmoid_table_225_3_sva | (~ initialized_sva);
  assign sigmoid_table_226_3_sva_dfm_1 = sigmoid_table_226_3_sva | (~ initialized_sva);
  assign sigmoid_table_227_3_sva_dfm_1 = sigmoid_table_227_3_sva | (~ initialized_sva);
  assign sigmoid_table_228_3_sva_dfm_1 = sigmoid_table_228_3_sva | (~ initialized_sva);
  assign sigmoid_table_274_3_sva_dfm_1 = sigmoid_table_274_3_sva | (~ initialized_sva);
  assign sigmoid_table_275_3_sva_dfm_1 = sigmoid_table_275_3_sva | (~ initialized_sva);
  assign sigmoid_table_276_3_sva_dfm_1 = sigmoid_table_276_3_sva | (~ initialized_sva);
  assign sigmoid_table_277_3_sva_dfm_1 = sigmoid_table_277_3_sva | (~ initialized_sva);
  assign sigmoid_table_278_3_sva_dfm_1 = sigmoid_table_278_3_sva | (~ initialized_sva);
  assign sigmoid_table_279_3_sva_dfm_1 = sigmoid_table_279_3_sva | (~ initialized_sva);
  assign sigmoid_table_280_3_sva_dfm_1 = sigmoid_table_280_3_sva | (~ initialized_sva);
  assign sigmoid_table_281_3_sva_dfm_1 = sigmoid_table_281_3_sva | (~ initialized_sva);
  assign sigmoid_table_282_3_sva_dfm_1 = sigmoid_table_282_3_sva | (~ initialized_sva);
  assign sigmoid_table_283_3_sva_dfm_1 = sigmoid_table_283_3_sva | (~ initialized_sva);
  assign sigmoid_table_308_3_sva_dfm_1 = sigmoid_table_308_3_sva | (~ initialized_sva);
  assign sigmoid_table_309_3_sva_dfm_1 = sigmoid_table_309_3_sva | (~ initialized_sva);
  assign sigmoid_table_310_3_sva_dfm_1 = sigmoid_table_310_3_sva | (~ initialized_sva);
  assign sigmoid_table_311_3_sva_dfm_1 = sigmoid_table_311_3_sva | (~ initialized_sva);
  assign sigmoid_table_312_3_sva_dfm_1 = sigmoid_table_312_3_sva | (~ initialized_sva);
  assign sigmoid_table_313_3_sva_dfm_1 = sigmoid_table_313_3_sva | (~ initialized_sva);
  assign sigmoid_table_330_3_sva_dfm_1 = sigmoid_table_330_3_sva | (~ initialized_sva);
  assign sigmoid_table_331_3_sva_dfm_1 = sigmoid_table_331_3_sva | (~ initialized_sva);
  assign sigmoid_table_332_3_sva_dfm_1 = sigmoid_table_332_3_sva | (~ initialized_sva);
  assign sigmoid_table_333_3_sva_dfm_1 = sigmoid_table_333_3_sva | (~ initialized_sva);
  assign sigmoid_table_334_3_sva_dfm_1 = sigmoid_table_334_3_sva | (~ initialized_sva);
  assign sigmoid_table_347_3_sva_dfm_1 = sigmoid_table_347_3_sva | (~ initialized_sva);
  assign sigmoid_table_348_3_sva_dfm_1 = sigmoid_table_348_3_sva | (~ initialized_sva);
  assign sigmoid_table_349_3_sva_dfm_1 = sigmoid_table_349_3_sva | (~ initialized_sva);
  assign sigmoid_table_350_3_sva_dfm_1 = sigmoid_table_350_3_sva | (~ initialized_sva);
  assign sigmoid_table_361_3_sva_dfm_1 = sigmoid_table_361_3_sva | (~ initialized_sva);
  assign sigmoid_table_362_3_sva_dfm_1 = sigmoid_table_362_3_sva | (~ initialized_sva);
  assign sigmoid_table_363_3_sva_dfm_1 = sigmoid_table_363_3_sva | (~ initialized_sva);
  assign sigmoid_table_373_3_sva_dfm_1 = sigmoid_table_373_3_sva | (~ initialized_sva);
  assign sigmoid_table_374_3_sva_dfm_1 = sigmoid_table_374_3_sva | (~ initialized_sva);
  assign sigmoid_table_375_3_sva_dfm_1 = sigmoid_table_375_3_sva | (~ initialized_sva);
  assign sigmoid_table_383_3_sva_dfm_1 = sigmoid_table_383_3_sva | (~ initialized_sva);
  assign sigmoid_table_384_3_sva_dfm_1 = sigmoid_table_384_3_sva | (~ initialized_sva);
  assign sigmoid_table_385_3_sva_dfm_1 = sigmoid_table_385_3_sva | (~ initialized_sva);
  assign sigmoid_table_392_3_sva_dfm_1 = sigmoid_table_392_3_sva | (~ initialized_sva);
  assign sigmoid_table_393_3_sva_dfm_1 = sigmoid_table_393_3_sva | (~ initialized_sva);
  assign sigmoid_table_394_3_sva_dfm_1 = sigmoid_table_394_3_sva | (~ initialized_sva);
  assign sigmoid_table_401_3_sva_dfm_1 = sigmoid_table_401_3_sva | (~ initialized_sva);
  assign sigmoid_table_402_3_sva_dfm_1 = sigmoid_table_402_3_sva | (~ initialized_sva);
  assign sigmoid_table_408_3_sva_dfm_1 = sigmoid_table_408_3_sva | (~ initialized_sva);
  assign sigmoid_table_409_3_sva_dfm_1 = sigmoid_table_409_3_sva | (~ initialized_sva);
  assign sigmoid_table_415_3_sva_dfm_1 = sigmoid_table_415_3_sva | (~ initialized_sva);
  assign sigmoid_table_416_3_sva_dfm_1 = sigmoid_table_416_3_sva | (~ initialized_sva);
  assign sigmoid_table_422_3_sva_dfm_1 = sigmoid_table_422_3_sva | (~ initialized_sva);
  assign sigmoid_table_428_3_sva_dfm_1 = sigmoid_table_428_3_sva | (~ initialized_sva);
  assign sigmoid_table_429_3_sva_dfm_1 = sigmoid_table_429_3_sva | (~ initialized_sva);
  assign sigmoid_table_434_3_sva_dfm_1 = sigmoid_table_434_3_sva | (~ initialized_sva);
  assign sigmoid_table_445_3_sva_dfm_1 = sigmoid_table_445_3_sva | (~ initialized_sva);
  assign sigmoid_table_450_3_sva_dfm_1 = sigmoid_table_450_3_sva | (~ initialized_sva);
  assign sigmoid_table_455_3_sva_dfm_1 = sigmoid_table_455_3_sva | (~ initialized_sva);
  assign sigmoid_table_460_3_sva_dfm_1 = sigmoid_table_460_3_sva | (~ initialized_sva);
  assign sigmoid_table_464_3_sva_dfm_1 = sigmoid_table_464_3_sva | (~ initialized_sva);
  assign sigmoid_table_469_3_sva_dfm_1 = sigmoid_table_469_3_sva | (~ initialized_sva);
  assign sigmoid_table_473_3_sva_dfm_1 = sigmoid_table_473_3_sva | (~ initialized_sva);
  assign sigmoid_table_478_3_sva_dfm_1 = sigmoid_table_478_3_sva | (~ initialized_sva);
  assign sigmoid_table_482_3_sva_dfm_1 = sigmoid_table_482_3_sva | (~ initialized_sva);
  assign sigmoid_table_486_3_sva_dfm_1 = sigmoid_table_486_3_sva | (~ initialized_sva);
  assign sigmoid_table_490_3_sva_dfm_1 = sigmoid_table_490_3_sva | (~ initialized_sva);
  assign sigmoid_table_494_3_sva_dfm_1 = sigmoid_table_494_3_sva | (~ initialized_sva);
  assign sigmoid_table_498_3_sva_dfm_1 = sigmoid_table_498_3_sva | (~ initialized_sva);
  assign sigmoid_table_502_3_sva_dfm_1 = sigmoid_table_502_3_sva | (~ initialized_sva);
  assign sigmoid_table_506_3_sva_dfm_1 = sigmoid_table_506_3_sva | (~ initialized_sva);
  assign sigmoid_table_514_3_sva_dfm_1 = sigmoid_table_514_3_sva | (~ initialized_sva);
  assign sigmoid_table_519_3_sva_dfm_1 = sigmoid_table_519_3_sva | (~ initialized_sva);
  assign sigmoid_table_523_3_sva_dfm_1 = sigmoid_table_523_3_sva | (~ initialized_sva);
  assign sigmoid_table_527_3_sva_dfm_1 = sigmoid_table_527_3_sva | (~ initialized_sva);
  assign sigmoid_table_531_3_sva_dfm_1 = sigmoid_table_531_3_sva | (~ initialized_sva);
  assign sigmoid_table_535_3_sva_dfm_1 = sigmoid_table_535_3_sva | (~ initialized_sva);
  assign sigmoid_table_539_3_sva_dfm_1 = sigmoid_table_539_3_sva | (~ initialized_sva);
  assign sigmoid_table_543_3_sva_dfm_1 = sigmoid_table_543_3_sva | (~ initialized_sva);
  assign sigmoid_table_547_3_sva_dfm_1 = sigmoid_table_547_3_sva | (~ initialized_sva);
  assign sigmoid_table_552_3_sva_dfm_1 = sigmoid_table_552_3_sva | (~ initialized_sva);
  assign sigmoid_table_556_3_sva_dfm_1 = sigmoid_table_556_3_sva | (~ initialized_sva);
  assign sigmoid_table_561_3_sva_dfm_1 = sigmoid_table_561_3_sva | (~ initialized_sva);
  assign sigmoid_table_565_3_sva_dfm_1 = sigmoid_table_565_3_sva | (~ initialized_sva);
  assign sigmoid_table_570_3_sva_dfm_1 = sigmoid_table_570_3_sva | (~ initialized_sva);
  assign sigmoid_table_575_3_sva_dfm_1 = sigmoid_table_575_3_sva | (~ initialized_sva);
  assign sigmoid_table_586_3_sva_dfm_1 = sigmoid_table_586_3_sva | (~ initialized_sva);
  assign sigmoid_table_591_3_sva_dfm_1 = sigmoid_table_591_3_sva | (~ initialized_sva);
  assign sigmoid_table_592_3_sva_dfm_1 = sigmoid_table_592_3_sva | (~ initialized_sva);
  assign sigmoid_table_597_3_sva_dfm_1 = sigmoid_table_597_3_sva | (~ initialized_sva);
  assign sigmoid_table_603_3_sva_dfm_1 = sigmoid_table_603_3_sva | (~ initialized_sva);
  assign sigmoid_table_604_3_sva_dfm_1 = sigmoid_table_604_3_sva | (~ initialized_sva);
  assign sigmoid_table_610_3_sva_dfm_1 = sigmoid_table_610_3_sva | (~ initialized_sva);
  assign sigmoid_table_617_3_sva_dfm_1 = sigmoid_table_617_3_sva | (~ initialized_sva);
  assign sigmoid_table_618_3_sva_dfm_1 = sigmoid_table_618_3_sva | (~ initialized_sva);
  assign sigmoid_table_624_3_sva_dfm_1 = sigmoid_table_624_3_sva | (~ initialized_sva);
  assign sigmoid_table_625_3_sva_dfm_1 = sigmoid_table_625_3_sva | (~ initialized_sva);
  assign sigmoid_table_633_3_sva_dfm_1 = sigmoid_table_633_3_sva | (~ initialized_sva);
  assign sigmoid_table_634_3_sva_dfm_1 = sigmoid_table_634_3_sva | (~ initialized_sva);
  assign sigmoid_table_642_3_sva_dfm_1 = sigmoid_table_642_3_sva | (~ initialized_sva);
  assign sigmoid_table_643_3_sva_dfm_1 = sigmoid_table_643_3_sva | (~ initialized_sva);
  assign sigmoid_table_652_3_sva_dfm_1 = sigmoid_table_652_3_sva | (~ initialized_sva);
  assign sigmoid_table_653_3_sva_dfm_1 = sigmoid_table_653_3_sva | (~ initialized_sva);
  assign sigmoid_table_654_3_sva_dfm_1 = sigmoid_table_654_3_sva | (~ initialized_sva);
  assign sigmoid_table_664_3_sva_dfm_1 = sigmoid_table_664_3_sva | (~ initialized_sva);
  assign sigmoid_table_665_3_sva_dfm_1 = sigmoid_table_665_3_sva | (~ initialized_sva);
  assign sigmoid_table_666_3_sva_dfm_1 = sigmoid_table_666_3_sva | (~ initialized_sva);
  assign sigmoid_table_678_3_sva_dfm_1 = sigmoid_table_678_3_sva | (~ initialized_sva);
  assign sigmoid_table_679_3_sva_dfm_1 = sigmoid_table_679_3_sva | (~ initialized_sva);
  assign sigmoid_table_680_3_sva_dfm_1 = sigmoid_table_680_3_sva | (~ initialized_sva);
  assign sigmoid_table_681_3_sva_dfm_1 = sigmoid_table_681_3_sva | (~ initialized_sva);
  assign sigmoid_table_695_3_sva_dfm_1 = sigmoid_table_695_3_sva | (~ initialized_sva);
  assign sigmoid_table_696_3_sva_dfm_1 = sigmoid_table_696_3_sva | (~ initialized_sva);
  assign sigmoid_table_697_3_sva_dfm_1 = sigmoid_table_697_3_sva | (~ initialized_sva);
  assign sigmoid_table_698_3_sva_dfm_1 = sigmoid_table_698_3_sva | (~ initialized_sva);
  assign sigmoid_table_699_3_sva_dfm_1 = sigmoid_table_699_3_sva | (~ initialized_sva);
  assign sigmoid_table_717_3_sva_dfm_1 = sigmoid_table_717_3_sva | (~ initialized_sva);
  assign sigmoid_table_718_3_sva_dfm_1 = sigmoid_table_718_3_sva | (~ initialized_sva);
  assign sigmoid_table_719_3_sva_dfm_1 = sigmoid_table_719_3_sva | (~ initialized_sva);
  assign sigmoid_table_720_3_sva_dfm_1 = sigmoid_table_720_3_sva | (~ initialized_sva);
  assign sigmoid_table_721_3_sva_dfm_1 = sigmoid_table_721_3_sva | (~ initialized_sva);
  assign sigmoid_table_722_3_sva_dfm_1 = sigmoid_table_722_3_sva | (~ initialized_sva);
  assign sigmoid_table_723_3_sva_dfm_1 = sigmoid_table_723_3_sva | (~ initialized_sva);
  assign sigmoid_table_751_3_sva_dfm_1 = sigmoid_table_751_3_sva | (~ initialized_sva);
  assign sigmoid_table_752_3_sva_dfm_1 = sigmoid_table_752_3_sva | (~ initialized_sva);
  assign sigmoid_table_753_3_sva_dfm_1 = sigmoid_table_753_3_sva | (~ initialized_sva);
  assign sigmoid_table_754_3_sva_dfm_1 = sigmoid_table_754_3_sva | (~ initialized_sva);
  assign sigmoid_table_755_3_sva_dfm_1 = sigmoid_table_755_3_sva | (~ initialized_sva);
  assign sigmoid_table_756_3_sva_dfm_1 = sigmoid_table_756_3_sva | (~ initialized_sva);
  assign sigmoid_table_757_3_sva_dfm_1 = sigmoid_table_757_3_sva | (~ initialized_sva);
  assign sigmoid_table_758_3_sva_dfm_1 = sigmoid_table_758_3_sva | (~ initialized_sva);
  assign sigmoid_table_759_3_sva_dfm_1 = sigmoid_table_759_3_sva | (~ initialized_sva);
  assign sigmoid_table_760_3_sva_dfm_1 = sigmoid_table_760_3_sva | (~ initialized_sva);
  assign sigmoid_table_761_3_sva_dfm_1 = sigmoid_table_761_3_sva | (~ initialized_sva);
  assign sigmoid_table_762_3_sva_dfm_1 = sigmoid_table_762_3_sva | (~ initialized_sva);
  assign sigmoid_table_339_6_sva_dfm_1 = sigmoid_table_339_6_sva | (~ initialized_sva);
  assign sigmoid_table_340_6_sva_dfm_1 = sigmoid_table_340_6_sva | (~ initialized_sva);
  assign sigmoid_table_341_6_sva_dfm_1 = sigmoid_table_341_6_sva | (~ initialized_sva);
  assign sigmoid_table_342_6_sva_dfm_1 = sigmoid_table_342_6_sva | (~ initialized_sva);
  assign sigmoid_table_343_6_sva_dfm_1 = sigmoid_table_343_6_sva | (~ initialized_sva);
  assign sigmoid_table_344_6_sva_dfm_1 = sigmoid_table_344_6_sva | (~ initialized_sva);
  assign sigmoid_table_345_6_sva_dfm_1 = sigmoid_table_345_6_sva | (~ initialized_sva);
  assign sigmoid_table_346_6_sva_dfm_1 = sigmoid_table_346_6_sva | (~ initialized_sva);
  assign sigmoid_table_347_6_sva_dfm_1 = sigmoid_table_347_6_sva | (~ initialized_sva);
  assign sigmoid_table_348_6_sva_dfm_1 = sigmoid_table_348_6_sva | (~ initialized_sva);
  assign sigmoid_table_349_6_sva_dfm_1 = sigmoid_table_349_6_sva | (~ initialized_sva);
  assign sigmoid_table_350_6_sva_dfm_1 = sigmoid_table_350_6_sva | (~ initialized_sva);
  assign sigmoid_table_351_6_sva_dfm_1 = sigmoid_table_351_6_sva | (~ initialized_sva);
  assign sigmoid_table_352_6_sva_dfm_1 = sigmoid_table_352_6_sva | (~ initialized_sva);
  assign sigmoid_table_353_6_sva_dfm_1 = sigmoid_table_353_6_sva | (~ initialized_sva);
  assign sigmoid_table_354_6_sva_dfm_1 = sigmoid_table_354_6_sva | (~ initialized_sva);
  assign sigmoid_table_355_6_sva_dfm_1 = sigmoid_table_355_6_sva | (~ initialized_sva);
  assign sigmoid_table_356_6_sva_dfm_1 = sigmoid_table_356_6_sva | (~ initialized_sva);
  assign sigmoid_table_357_6_sva_dfm_1 = sigmoid_table_357_6_sva | (~ initialized_sva);
  assign sigmoid_table_358_6_sva_dfm_1 = sigmoid_table_358_6_sva | (~ initialized_sva);
  assign sigmoid_table_359_6_sva_dfm_1 = sigmoid_table_359_6_sva | (~ initialized_sva);
  assign sigmoid_table_360_6_sva_dfm_1 = sigmoid_table_360_6_sva | (~ initialized_sva);
  assign sigmoid_table_361_6_sva_dfm_1 = sigmoid_table_361_6_sva | (~ initialized_sva);
  assign sigmoid_table_362_6_sva_dfm_1 = sigmoid_table_362_6_sva | (~ initialized_sva);
  assign sigmoid_table_363_6_sva_dfm_1 = sigmoid_table_363_6_sva | (~ initialized_sva);
  assign sigmoid_table_364_6_sva_dfm_1 = sigmoid_table_364_6_sva | (~ initialized_sva);
  assign sigmoid_table_365_6_sva_dfm_1 = sigmoid_table_365_6_sva | (~ initialized_sva);
  assign sigmoid_table_366_6_sva_dfm_1 = sigmoid_table_366_6_sva | (~ initialized_sva);
  assign sigmoid_table_367_5_sva_dfm_1 = sigmoid_table_367_5_sva | (~ initialized_sva);
  assign sigmoid_table_368_5_sva_dfm_1 = sigmoid_table_368_5_sva | (~ initialized_sva);
  assign sigmoid_table_369_5_sva_dfm_1 = sigmoid_table_369_5_sva | (~ initialized_sva);
  assign sigmoid_table_370_5_sva_dfm_1 = sigmoid_table_370_5_sva | (~ initialized_sva);
  assign sigmoid_table_371_5_sva_dfm_1 = sigmoid_table_371_5_sva | (~ initialized_sva);
  assign sigmoid_table_372_5_sva_dfm_1 = sigmoid_table_372_5_sva | (~ initialized_sva);
  assign sigmoid_table_373_5_sva_dfm_1 = sigmoid_table_373_5_sva | (~ initialized_sva);
  assign sigmoid_table_374_5_sva_dfm_1 = sigmoid_table_374_5_sva | (~ initialized_sva);
  assign sigmoid_table_375_5_sva_dfm_1 = sigmoid_table_375_5_sva | (~ initialized_sva);
  assign sigmoid_table_376_5_sva_dfm_1 = sigmoid_table_376_5_sva | (~ initialized_sva);
  assign sigmoid_table_377_5_sva_dfm_1 = sigmoid_table_377_5_sva | (~ initialized_sva);
  assign sigmoid_table_378_4_sva_dfm_1 = sigmoid_table_378_4_sva | (~ initialized_sva);
  assign sigmoid_table_379_4_sva_dfm_1 = sigmoid_table_379_4_sva | (~ initialized_sva);
  assign sigmoid_table_380_4_sva_dfm_1 = sigmoid_table_380_4_sva | (~ initialized_sva);
  assign sigmoid_table_381_4_sva_dfm_1 = sigmoid_table_381_4_sva | (~ initialized_sva);
  assign sigmoid_table_382_4_sva_dfm_1 = sigmoid_table_382_4_sva | (~ initialized_sva);
  assign sigmoid_table_462_6_sva_dfm_1 = sigmoid_table_462_6_sva | (~ initialized_sva);
  assign sigmoid_table_463_6_sva_dfm_1 = sigmoid_table_463_6_sva | (~ initialized_sva);
  assign sigmoid_table_464_6_sva_dfm_1 = sigmoid_table_464_6_sva | (~ initialized_sva);
  assign sigmoid_table_465_6_sva_dfm_1 = sigmoid_table_465_6_sva | (~ initialized_sva);
  assign sigmoid_table_466_6_sva_dfm_1 = sigmoid_table_466_6_sva | (~ initialized_sva);
  assign sigmoid_table_467_6_sva_dfm_1 = sigmoid_table_467_6_sva | (~ initialized_sva);
  assign sigmoid_table_468_6_sva_dfm_1 = sigmoid_table_468_6_sva | (~ initialized_sva);
  assign sigmoid_table_469_6_sva_dfm_1 = sigmoid_table_469_6_sva | (~ initialized_sva);
  assign sigmoid_table_470_6_sva_dfm_1 = sigmoid_table_470_6_sva | (~ initialized_sva);
  assign sigmoid_table_471_5_sva_dfm_1 = sigmoid_table_471_5_sva | (~ initialized_sva);
  assign sigmoid_table_472_5_sva_dfm_1 = sigmoid_table_472_5_sva | (~ initialized_sva);
  assign sigmoid_table_473_5_sva_dfm_1 = sigmoid_table_473_5_sva | (~ initialized_sva);
  assign sigmoid_table_474_5_sva_dfm_1 = sigmoid_table_474_5_sva | (~ initialized_sva);
  assign sigmoid_table_475_5_sva_dfm_1 = sigmoid_table_475_5_sva | (~ initialized_sva);
  assign sigmoid_table_476_4_sva_dfm_1 = sigmoid_table_476_4_sva | (~ initialized_sva);
  assign sigmoid_table_477_4_sva_dfm_1 = sigmoid_table_477_4_sva | (~ initialized_sva);
  assign sigmoid_table_529_6_sva_dfm_1 = sigmoid_table_529_6_sva | (~ initialized_sva);
  assign sigmoid_table_530_6_sva_dfm_1 = sigmoid_table_530_6_sva | (~ initialized_sva);
  assign sigmoid_table_531_6_sva_dfm_1 = sigmoid_table_531_6_sva | (~ initialized_sva);
  assign sigmoid_table_532_6_sva_dfm_1 = sigmoid_table_532_6_sva | (~ initialized_sva);
  assign sigmoid_table_533_6_sva_dfm_1 = sigmoid_table_533_6_sva | (~ initialized_sva);
  assign sigmoid_table_534_6_sva_dfm_1 = sigmoid_table_534_6_sva | (~ initialized_sva);
  assign sigmoid_table_535_6_sva_dfm_1 = sigmoid_table_535_6_sva | (~ initialized_sva);
  assign sigmoid_table_536_6_sva_dfm_1 = sigmoid_table_536_6_sva | (~ initialized_sva);
  assign sigmoid_table_537_5_sva_dfm_1 = sigmoid_table_537_5_sva | (~ initialized_sva);
  assign sigmoid_table_538_5_sva_dfm_1 = sigmoid_table_538_5_sva | (~ initialized_sva);
  assign sigmoid_table_539_5_sva_dfm_1 = sigmoid_table_539_5_sva | (~ initialized_sva);
  assign sigmoid_table_540_5_sva_dfm_1 = sigmoid_table_540_5_sva | (~ initialized_sva);
  assign sigmoid_table_541_4_sva_dfm_1 = sigmoid_table_541_4_sva | (~ initialized_sva);
  assign sigmoid_table_542_4_sva_dfm_1 = sigmoid_table_542_4_sva | (~ initialized_sva);
  assign sigmoid_table_606_6_sva_dfm_1 = sigmoid_table_606_6_sva | (~ initialized_sva);
  assign sigmoid_table_607_6_sva_dfm_1 = sigmoid_table_607_6_sva | (~ initialized_sva);
  assign sigmoid_table_608_6_sva_dfm_1 = sigmoid_table_608_6_sva | (~ initialized_sva);
  assign sigmoid_table_609_6_sva_dfm_1 = sigmoid_table_609_6_sva | (~ initialized_sva);
  assign sigmoid_table_610_6_sva_dfm_1 = sigmoid_table_610_6_sva | (~ initialized_sva);
  assign sigmoid_table_611_6_sva_dfm_1 = sigmoid_table_611_6_sva | (~ initialized_sva);
  assign sigmoid_table_612_6_sva_dfm_1 = sigmoid_table_612_6_sva | (~ initialized_sva);
  assign sigmoid_table_613_6_sva_dfm_1 = sigmoid_table_613_6_sva | (~ initialized_sva);
  assign sigmoid_table_614_6_sva_dfm_1 = sigmoid_table_614_6_sva | (~ initialized_sva);
  assign sigmoid_table_615_6_sva_dfm_1 = sigmoid_table_615_6_sva | (~ initialized_sva);
  assign sigmoid_table_616_6_sva_dfm_1 = sigmoid_table_616_6_sva | (~ initialized_sva);
  assign sigmoid_table_617_6_sva_dfm_1 = sigmoid_table_617_6_sva | (~ initialized_sva);
  assign sigmoid_table_618_6_sva_dfm_1 = sigmoid_table_618_6_sva | (~ initialized_sva);
  assign sigmoid_table_619_6_sva_dfm_1 = sigmoid_table_619_6_sva | (~ initialized_sva);
  assign sigmoid_table_620_5_sva_dfm_1 = sigmoid_table_620_5_sva | (~ initialized_sva);
  assign sigmoid_table_621_5_sva_dfm_1 = sigmoid_table_621_5_sva | (~ initialized_sva);
  assign sigmoid_table_622_5_sva_dfm_1 = sigmoid_table_622_5_sva | (~ initialized_sva);
  assign sigmoid_table_623_5_sva_dfm_1 = sigmoid_table_623_5_sva | (~ initialized_sva);
  assign sigmoid_table_624_5_sva_dfm_1 = sigmoid_table_624_5_sva | (~ initialized_sva);
  assign sigmoid_table_625_5_sva_dfm_1 = sigmoid_table_625_5_sva | (~ initialized_sva);
  assign sigmoid_table_626_5_sva_dfm_1 = sigmoid_table_626_5_sva | (~ initialized_sva);
  assign sigmoid_table_627_5_sva_dfm_1 = sigmoid_table_627_5_sva | (~ initialized_sva);
  assign sigmoid_table_628_4_sva_dfm_1 = sigmoid_table_628_4_sva | (~ initialized_sva);
  assign sigmoid_table_629_4_sva_dfm_1 = sigmoid_table_629_4_sva | (~ initialized_sva);
  assign sigmoid_table_630_4_sva_dfm_1 = sigmoid_table_630_4_sva | (~ initialized_sva);
  assign sigmoid_table_631_4_sva_dfm_1 = sigmoid_table_631_4_sva | (~ initialized_sva);
  assign sigmoid_table_632_4_sva_dfm_1 = sigmoid_table_632_4_sva | (~ initialized_sva);
  assign sigmoid_table_247_4_sva_dfm_1 = sigmoid_table_247_4_sva | (~ initialized_sva);
  assign sigmoid_table_248_4_sva_dfm_1 = sigmoid_table_248_4_sva | (~ initialized_sva);
  assign sigmoid_table_249_4_sva_dfm_1 = sigmoid_table_249_4_sva | (~ initialized_sva);
  assign sigmoid_table_250_4_sva_dfm_1 = sigmoid_table_250_4_sva | (~ initialized_sva);
  assign sigmoid_table_251_4_sva_dfm_1 = sigmoid_table_251_4_sva | (~ initialized_sva);
  assign sigmoid_table_252_4_sva_dfm_1 = sigmoid_table_252_4_sva | (~ initialized_sva);
  assign sigmoid_table_253_4_sva_dfm_1 = sigmoid_table_253_4_sva | (~ initialized_sva);
  assign sigmoid_table_254_4_sva_dfm_1 = sigmoid_table_254_4_sva | (~ initialized_sva);
  assign sigmoid_table_255_4_sva_dfm_1 = sigmoid_table_255_4_sva | (~ initialized_sva);
  assign sigmoid_table_256_4_sva_dfm_1 = sigmoid_table_256_4_sva | (~ initialized_sva);
  assign sigmoid_table_257_4_sva_dfm_1 = sigmoid_table_257_4_sva | (~ initialized_sva);
  assign sigmoid_table_258_4_sva_dfm_1 = sigmoid_table_258_4_sva | (~ initialized_sva);
  assign sigmoid_table_259_4_sva_dfm_1 = sigmoid_table_259_4_sva | (~ initialized_sva);
  assign sigmoid_table_260_4_sva_dfm_1 = sigmoid_table_260_4_sva | (~ initialized_sva);
  assign sigmoid_table_261_4_sva_dfm_1 = sigmoid_table_261_4_sva | (~ initialized_sva);
  assign sigmoid_table_262_4_sva_dfm_1 = sigmoid_table_262_4_sva | (~ initialized_sva);
  assign sigmoid_table_263_4_sva_dfm_1 = sigmoid_table_263_4_sva | (~ initialized_sva);
  assign sigmoid_table_264_4_sva_dfm_1 = sigmoid_table_264_4_sva | (~ initialized_sva);
  assign sigmoid_table_265_4_sva_dfm_1 = sigmoid_table_265_4_sva | (~ initialized_sva);
  assign sigmoid_table_266_4_sva_dfm_1 = sigmoid_table_266_4_sva | (~ initialized_sva);
  assign sigmoid_table_267_4_sva_dfm_1 = sigmoid_table_267_4_sva | (~ initialized_sva);
  assign sigmoid_table_268_4_sva_dfm_1 = sigmoid_table_268_4_sva | (~ initialized_sva);
  assign sigmoid_table_269_4_sva_dfm_1 = sigmoid_table_269_4_sva | (~ initialized_sva);
  assign sigmoid_table_270_4_sva_dfm_1 = sigmoid_table_270_4_sva | (~ initialized_sva);
  assign sigmoid_table_271_4_sva_dfm_1 = sigmoid_table_271_4_sva | (~ initialized_sva);
  assign sigmoid_table_272_4_sva_dfm_1 = sigmoid_table_272_4_sva | (~ initialized_sva);
  assign sigmoid_table_273_4_sva_dfm_1 = sigmoid_table_273_4_sva | (~ initialized_sva);
  assign sigmoid_table_320_4_sva_dfm_1 = sigmoid_table_320_4_sva | (~ initialized_sva);
  assign sigmoid_table_321_4_sva_dfm_1 = sigmoid_table_321_4_sva | (~ initialized_sva);
  assign sigmoid_table_322_4_sva_dfm_1 = sigmoid_table_322_4_sva | (~ initialized_sva);
  assign sigmoid_table_323_4_sva_dfm_1 = sigmoid_table_323_4_sva | (~ initialized_sva);
  assign sigmoid_table_324_4_sva_dfm_1 = sigmoid_table_324_4_sva | (~ initialized_sva);
  assign sigmoid_table_325_4_sva_dfm_1 = sigmoid_table_325_4_sva | (~ initialized_sva);
  assign sigmoid_table_326_4_sva_dfm_1 = sigmoid_table_326_4_sva | (~ initialized_sva);
  assign sigmoid_table_327_4_sva_dfm_1 = sigmoid_table_327_4_sva | (~ initialized_sva);
  assign sigmoid_table_328_4_sva_dfm_1 = sigmoid_table_328_4_sva | (~ initialized_sva);
  assign sigmoid_table_329_4_sva_dfm_1 = sigmoid_table_329_4_sva | (~ initialized_sva);
  assign sigmoid_table_355_4_sva_dfm_1 = sigmoid_table_355_4_sva | (~ initialized_sva);
  assign sigmoid_table_356_4_sva_dfm_1 = sigmoid_table_356_4_sva | (~ initialized_sva);
  assign sigmoid_table_357_4_sva_dfm_1 = sigmoid_table_357_4_sva | (~ initialized_sva);
  assign sigmoid_table_358_4_sva_dfm_1 = sigmoid_table_358_4_sva | (~ initialized_sva);
  assign sigmoid_table_359_4_sva_dfm_1 = sigmoid_table_359_4_sva | (~ initialized_sva);
  assign sigmoid_table_360_4_sva_dfm_1 = sigmoid_table_360_4_sva | (~ initialized_sva);
  assign sigmoid_table_397_4_sva_dfm_1 = sigmoid_table_397_4_sva | (~ initialized_sva);
  assign sigmoid_table_398_4_sva_dfm_1 = sigmoid_table_398_4_sva | (~ initialized_sva);
  assign sigmoid_table_399_4_sva_dfm_1 = sigmoid_table_399_4_sva | (~ initialized_sva);
  assign sigmoid_table_400_4_sva_dfm_1 = sigmoid_table_400_4_sva | (~ initialized_sva);
  assign sigmoid_table_412_4_sva_dfm_1 = sigmoid_table_412_4_sva | (~ initialized_sva);
  assign sigmoid_table_413_4_sva_dfm_1 = sigmoid_table_413_4_sva | (~ initialized_sva);
  assign sigmoid_table_414_4_sva_dfm_1 = sigmoid_table_414_4_sva | (~ initialized_sva);
  assign sigmoid_table_425_4_sva_dfm_1 = sigmoid_table_425_4_sva | (~ initialized_sva);
  assign sigmoid_table_426_4_sva_dfm_1 = sigmoid_table_426_4_sva | (~ initialized_sva);
  assign sigmoid_table_427_4_sva_dfm_1 = sigmoid_table_427_4_sva | (~ initialized_sva);
  assign sigmoid_table_447_4_sva_dfm_1 = sigmoid_table_447_4_sva | (~ initialized_sva);
  assign sigmoid_table_448_4_sva_dfm_1 = sigmoid_table_448_4_sva | (~ initialized_sva);
  assign sigmoid_table_449_4_sva_dfm_1 = sigmoid_table_449_4_sva | (~ initialized_sva);
  assign sigmoid_table_457_4_sva_dfm_1 = sigmoid_table_457_4_sva | (~ initialized_sva);
  assign sigmoid_table_458_4_sva_dfm_1 = sigmoid_table_458_4_sva | (~ initialized_sva);
  assign sigmoid_table_459_4_sva_dfm_1 = sigmoid_table_459_4_sva | (~ initialized_sva);
  assign sigmoid_table_467_4_sva_dfm_1 = sigmoid_table_467_4_sva | (~ initialized_sva);
  assign sigmoid_table_468_4_sva_dfm_1 = sigmoid_table_468_4_sva | (~ initialized_sva);
  assign sigmoid_table_484_4_sva_dfm_1 = sigmoid_table_484_4_sva | (~ initialized_sva);
  assign sigmoid_table_485_4_sva_dfm_1 = sigmoid_table_485_4_sva | (~ initialized_sva);
  assign sigmoid_table_492_4_sva_dfm_1 = sigmoid_table_492_4_sva | (~ initialized_sva);
  assign sigmoid_table_493_4_sva_dfm_1 = sigmoid_table_493_4_sva | (~ initialized_sva);
  assign sigmoid_table_500_4_sva_dfm_1 = sigmoid_table_500_4_sva | (~ initialized_sva);
  assign sigmoid_table_501_4_sva_dfm_1 = sigmoid_table_501_4_sva | (~ initialized_sva);
  assign sigmoid_table_517_4_sva_dfm_1 = sigmoid_table_517_4_sva | (~ initialized_sva);
  assign sigmoid_table_518_4_sva_dfm_1 = sigmoid_table_518_4_sva | (~ initialized_sva);
  assign sigmoid_table_525_4_sva_dfm_1 = sigmoid_table_525_4_sva | (~ initialized_sva);
  assign sigmoid_table_526_4_sva_dfm_1 = sigmoid_table_526_4_sva | (~ initialized_sva);
  assign sigmoid_table_533_4_sva_dfm_1 = sigmoid_table_533_4_sva | (~ initialized_sva);
  assign sigmoid_table_534_4_sva_dfm_1 = sigmoid_table_534_4_sva | (~ initialized_sva);
  assign sigmoid_table_549_4_sva_dfm_1 = sigmoid_table_549_4_sva | (~ initialized_sva);
  assign sigmoid_table_550_4_sva_dfm_1 = sigmoid_table_550_4_sva | (~ initialized_sva);
  assign sigmoid_table_551_4_sva_dfm_1 = sigmoid_table_551_4_sva | (~ initialized_sva);
  assign sigmoid_table_558_4_sva_dfm_1 = sigmoid_table_558_4_sva | (~ initialized_sva);
  assign sigmoid_table_559_4_sva_dfm_1 = sigmoid_table_559_4_sva | (~ initialized_sva);
  assign sigmoid_table_560_4_sva_dfm_1 = sigmoid_table_560_4_sva | (~ initialized_sva);
  assign sigmoid_table_568_4_sva_dfm_1 = sigmoid_table_568_4_sva | (~ initialized_sva);
  assign sigmoid_table_569_4_sva_dfm_1 = sigmoid_table_569_4_sva | (~ initialized_sva);
  assign sigmoid_table_588_4_sva_dfm_1 = sigmoid_table_588_4_sva | (~ initialized_sva);
  assign sigmoid_table_589_4_sva_dfm_1 = sigmoid_table_589_4_sva | (~ initialized_sva);
  assign sigmoid_table_590_4_sva_dfm_1 = sigmoid_table_590_4_sva | (~ initialized_sva);
  assign sigmoid_table_600_4_sva_dfm_1 = sigmoid_table_600_4_sva | (~ initialized_sva);
  assign sigmoid_table_601_4_sva_dfm_1 = sigmoid_table_601_4_sva | (~ initialized_sva);
  assign sigmoid_table_602_4_sva_dfm_1 = sigmoid_table_602_4_sva | (~ initialized_sva);
  assign sigmoid_table_613_4_sva_dfm_1 = sigmoid_table_613_4_sva | (~ initialized_sva);
  assign sigmoid_table_614_4_sva_dfm_1 = sigmoid_table_614_4_sva | (~ initialized_sva);
  assign sigmoid_table_615_4_sva_dfm_1 = sigmoid_table_615_4_sva | (~ initialized_sva);
  assign sigmoid_table_616_4_sva_dfm_1 = sigmoid_table_616_4_sva | (~ initialized_sva);
  assign sigmoid_table_647_4_sva_dfm_1 = sigmoid_table_647_4_sva | (~ initialized_sva);
  assign sigmoid_table_648_4_sva_dfm_1 = sigmoid_table_648_4_sva | (~ initialized_sva);
  assign sigmoid_table_649_4_sva_dfm_1 = sigmoid_table_649_4_sva | (~ initialized_sva);
  assign sigmoid_table_650_4_sva_dfm_1 = sigmoid_table_650_4_sva | (~ initialized_sva);
  assign sigmoid_table_651_4_sva_dfm_1 = sigmoid_table_651_4_sva | (~ initialized_sva);
  assign sigmoid_table_670_4_sva_dfm_1 = sigmoid_table_670_4_sva | (~ initialized_sva);
  assign sigmoid_table_671_4_sva_dfm_1 = sigmoid_table_671_4_sva | (~ initialized_sva);
  assign sigmoid_table_672_4_sva_dfm_1 = sigmoid_table_672_4_sva | (~ initialized_sva);
  assign sigmoid_table_673_4_sva_dfm_1 = sigmoid_table_673_4_sva | (~ initialized_sva);
  assign sigmoid_table_674_4_sva_dfm_1 = sigmoid_table_674_4_sva | (~ initialized_sva);
  assign sigmoid_table_675_4_sva_dfm_1 = sigmoid_table_675_4_sva | (~ initialized_sva);
  assign sigmoid_table_676_4_sva_dfm_1 = sigmoid_table_676_4_sva | (~ initialized_sva);
  assign sigmoid_table_677_4_sva_dfm_1 = sigmoid_table_677_4_sva | (~ initialized_sva);
  assign sigmoid_table_705_4_sva_dfm_1 = sigmoid_table_705_4_sva | (~ initialized_sva);
  assign sigmoid_table_706_4_sva_dfm_1 = sigmoid_table_706_4_sva | (~ initialized_sva);
  assign sigmoid_table_707_4_sva_dfm_1 = sigmoid_table_707_4_sva | (~ initialized_sva);
  assign sigmoid_table_708_4_sva_dfm_1 = sigmoid_table_708_4_sva | (~ initialized_sva);
  assign sigmoid_table_709_4_sva_dfm_1 = sigmoid_table_709_4_sva | (~ initialized_sva);
  assign sigmoid_table_710_4_sva_dfm_1 = sigmoid_table_710_4_sva | (~ initialized_sva);
  assign sigmoid_table_711_4_sva_dfm_1 = sigmoid_table_711_4_sva | (~ initialized_sva);
  assign sigmoid_table_712_4_sva_dfm_1 = sigmoid_table_712_4_sva | (~ initialized_sva);
  assign sigmoid_table_713_4_sva_dfm_1 = sigmoid_table_713_4_sva | (~ initialized_sva);
  assign sigmoid_table_714_4_sva_dfm_1 = sigmoid_table_714_4_sva | (~ initialized_sva);
  assign sigmoid_table_715_4_sva_dfm_1 = sigmoid_table_715_4_sva | (~ initialized_sva);
  assign sigmoid_table_716_4_sva_dfm_1 = sigmoid_table_716_4_sva | (~ initialized_sva);
  assign sigmoid_table_293_5_sva_dfm_1 = sigmoid_table_293_5_sva | (~ initialized_sva);
  assign sigmoid_table_294_5_sva_dfm_1 = sigmoid_table_294_5_sva | (~ initialized_sva);
  assign sigmoid_table_295_5_sva_dfm_1 = sigmoid_table_295_5_sva | (~ initialized_sva);
  assign sigmoid_table_296_5_sva_dfm_1 = sigmoid_table_296_5_sva | (~ initialized_sva);
  assign sigmoid_table_297_5_sva_dfm_1 = sigmoid_table_297_5_sva | (~ initialized_sva);
  assign sigmoid_table_298_5_sva_dfm_1 = sigmoid_table_298_5_sva | (~ initialized_sva);
  assign sigmoid_table_299_5_sva_dfm_1 = sigmoid_table_299_5_sva | (~ initialized_sva);
  assign sigmoid_table_300_5_sva_dfm_1 = sigmoid_table_300_5_sva | (~ initialized_sva);
  assign sigmoid_table_301_5_sva_dfm_1 = sigmoid_table_301_5_sva | (~ initialized_sva);
  assign sigmoid_table_302_5_sva_dfm_1 = sigmoid_table_302_5_sva | (~ initialized_sva);
  assign sigmoid_table_303_5_sva_dfm_1 = sigmoid_table_303_5_sva | (~ initialized_sva);
  assign sigmoid_table_304_5_sva_dfm_1 = sigmoid_table_304_5_sva | (~ initialized_sva);
  assign sigmoid_table_305_5_sva_dfm_1 = sigmoid_table_305_5_sva | (~ initialized_sva);
  assign sigmoid_table_306_5_sva_dfm_1 = sigmoid_table_306_5_sva | (~ initialized_sva);
  assign sigmoid_table_307_5_sva_dfm_1 = sigmoid_table_307_5_sva | (~ initialized_sva);
  assign sigmoid_table_308_5_sva_dfm_1 = sigmoid_table_308_5_sva | (~ initialized_sva);
  assign sigmoid_table_309_5_sva_dfm_1 = sigmoid_table_309_5_sva | (~ initialized_sva);
  assign sigmoid_table_310_5_sva_dfm_1 = sigmoid_table_310_5_sva | (~ initialized_sva);
  assign sigmoid_table_311_5_sva_dfm_1 = sigmoid_table_311_5_sva | (~ initialized_sva);
  assign sigmoid_table_312_5_sva_dfm_1 = sigmoid_table_312_5_sva | (~ initialized_sva);
  assign sigmoid_table_313_5_sva_dfm_1 = sigmoid_table_313_5_sva | (~ initialized_sva);
  assign sigmoid_table_314_5_sva_dfm_1 = sigmoid_table_314_5_sva | (~ initialized_sva);
  assign sigmoid_table_315_5_sva_dfm_1 = sigmoid_table_315_5_sva | (~ initialized_sva);
  assign sigmoid_table_316_5_sva_dfm_1 = sigmoid_table_316_5_sva | (~ initialized_sva);
  assign sigmoid_table_317_5_sva_dfm_1 = sigmoid_table_317_5_sva | (~ initialized_sva);
  assign sigmoid_table_318_5_sva_dfm_1 = sigmoid_table_318_5_sva | (~ initialized_sva);
  assign sigmoid_table_319_5_sva_dfm_1 = sigmoid_table_319_5_sva | (~ initialized_sva);
  assign sigmoid_table_405_5_sva_dfm_1 = sigmoid_table_405_5_sva | (~ initialized_sva);
  assign sigmoid_table_406_5_sva_dfm_1 = sigmoid_table_406_5_sva | (~ initialized_sva);
  assign sigmoid_table_407_5_sva_dfm_1 = sigmoid_table_407_5_sva | (~ initialized_sva);
  assign sigmoid_table_408_5_sva_dfm_1 = sigmoid_table_408_5_sva | (~ initialized_sva);
  assign sigmoid_table_409_5_sva_dfm_1 = sigmoid_table_409_5_sva | (~ initialized_sva);
  assign sigmoid_table_410_5_sva_dfm_1 = sigmoid_table_410_5_sva | (~ initialized_sva);
  assign sigmoid_table_411_5_sva_dfm_1 = sigmoid_table_411_5_sva | (~ initialized_sva);
  assign sigmoid_table_452_5_sva_dfm_1 = sigmoid_table_452_5_sva | (~ initialized_sva);
  assign sigmoid_table_453_5_sva_dfm_1 = sigmoid_table_453_5_sva | (~ initialized_sva);
  assign sigmoid_table_454_5_sva_dfm_1 = sigmoid_table_454_5_sva | (~ initialized_sva);
  assign sigmoid_table_455_5_sva_dfm_1 = sigmoid_table_455_5_sva | (~ initialized_sva);
  assign sigmoid_table_456_5_sva_dfm_1 = sigmoid_table_456_5_sva | (~ initialized_sva);
  assign sigmoid_table_488_5_sva_dfm_1 = sigmoid_table_488_5_sva | (~ initialized_sva);
  assign sigmoid_table_489_5_sva_dfm_1 = sigmoid_table_489_5_sva | (~ initialized_sva);
  assign sigmoid_table_490_5_sva_dfm_1 = sigmoid_table_490_5_sva | (~ initialized_sva);
  assign sigmoid_table_491_5_sva_dfm_1 = sigmoid_table_491_5_sva | (~ initialized_sva);
  assign sigmoid_table_521_5_sva_dfm_1 = sigmoid_table_521_5_sva | (~ initialized_sva);
  assign sigmoid_table_522_5_sva_dfm_1 = sigmoid_table_522_5_sva | (~ initialized_sva);
  assign sigmoid_table_523_5_sva_dfm_1 = sigmoid_table_523_5_sva | (~ initialized_sva);
  assign sigmoid_table_524_5_sva_dfm_1 = sigmoid_table_524_5_sva | (~ initialized_sva);
  assign sigmoid_table_554_5_sva_dfm_1 = sigmoid_table_554_5_sva | (~ initialized_sva);
  assign sigmoid_table_555_5_sva_dfm_1 = sigmoid_table_555_5_sva | (~ initialized_sva);
  assign sigmoid_table_556_5_sva_dfm_1 = sigmoid_table_556_5_sva | (~ initialized_sva);
  assign sigmoid_table_557_5_sva_dfm_1 = sigmoid_table_557_5_sva | (~ initialized_sva);
  assign sigmoid_table_594_5_sva_dfm_1 = sigmoid_table_594_5_sva | (~ initialized_sva);
  assign sigmoid_table_595_5_sva_dfm_1 = sigmoid_table_595_5_sva | (~ initialized_sva);
  assign sigmoid_table_596_5_sva_dfm_1 = sigmoid_table_596_5_sva | (~ initialized_sva);
  assign sigmoid_table_597_5_sva_dfm_1 = sigmoid_table_597_5_sva | (~ initialized_sva);
  assign sigmoid_table_598_5_sva_dfm_1 = sigmoid_table_598_5_sva | (~ initialized_sva);
  assign sigmoid_table_599_5_sva_dfm_1 = sigmoid_table_599_5_sva | (~ initialized_sva);
  assign sigmoid_table_658_5_sva_dfm_1 = sigmoid_table_658_5_sva | (~ initialized_sva);
  assign sigmoid_table_659_5_sva_dfm_1 = sigmoid_table_659_5_sva | (~ initialized_sva);
  assign sigmoid_table_660_5_sva_dfm_1 = sigmoid_table_660_5_sva | (~ initialized_sva);
  assign sigmoid_table_661_5_sva_dfm_1 = sigmoid_table_661_5_sva | (~ initialized_sva);
  assign sigmoid_table_662_5_sva_dfm_1 = sigmoid_table_662_5_sva | (~ initialized_sva);
  assign sigmoid_table_663_5_sva_dfm_1 = sigmoid_table_663_5_sva | (~ initialized_sva);
  assign sigmoid_table_664_5_sva_dfm_1 = sigmoid_table_664_5_sva | (~ initialized_sva);
  assign sigmoid_table_665_5_sva_dfm_1 = sigmoid_table_665_5_sva | (~ initialized_sva);
  assign sigmoid_table_666_5_sva_dfm_1 = sigmoid_table_666_5_sva | (~ initialized_sva);
  assign sigmoid_table_667_5_sva_dfm_1 = sigmoid_table_667_5_sva | (~ initialized_sva);
  assign sigmoid_table_668_5_sva_dfm_1 = sigmoid_table_668_5_sva | (~ initialized_sva);
  assign sigmoid_table_669_5_sva_dfm_1 = sigmoid_table_669_5_sva | (~ initialized_sva);
  assign nl_operator_32_true_acc_psp_sva_1 = conv_s2s_5_6(data_rsci_idat[17:13])
      + 6'b000001;
  assign operator_32_true_acc_psp_sva_1 = nl_operator_32_true_acc_psp_sva_1[5:0];
  assign nl_operator_32_true_acc_nl =  -(index_14_9_lpi_1_dfm_1[5:1]);
  assign operator_32_true_acc_nl = nl_operator_32_true_acc_nl[4:0];
  assign operator_32_true_acc_itm_4 = readslicef_5_1_4((operator_32_true_acc_nl));
  assign operator_32_true_not_2_nl = ~ (operator_32_true_acc_psp_sva_1[5]);
  assign index_14_9_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, operator_32_true_acc_psp_sva_1,
      (operator_32_true_not_2_nl));
  assign for_for_or_1_itm = (index_14_9_lpi_1_dfm_1[0]) | operator_32_true_acc_itm_4;
  assign operator_32_true_not_4_nl = ~ (operator_32_true_acc_psp_sva_1[5]);
  assign for_for_and_1_nl = MUX_v_9_2_2(9'b000000000, (data_rsci_idat[12:4]), (operator_32_true_not_4_nl));
  assign for_for_or_itm = MUX_v_9_2_2((for_for_and_1_nl), 9'b111111111, operator_32_true_acc_itm_4);
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      res_rsci_d_0 <= 1'b0;
      res_rsci_d_9 <= 1'b0;
      res_rsci_d_1 <= 1'b0;
      res_rsci_d_8 <= 1'b0;
      res_rsci_d_2 <= 1'b0;
      res_rsci_d_7 <= 1'b0;
      res_rsci_d_3 <= 1'b0;
      res_rsci_d_6 <= 1'b0;
      res_rsci_d_4 <= 1'b0;
      res_rsci_d_5 <= 1'b0;
      initialized_sva <= 1'b0;
    end
    else if ( ccs_ccore_en ) begin
      res_rsci_d_0 <= MUX_s_1_1024_2(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, sigmoid_table_69_0_sva_dfm_1, sigmoid_table_70_0_sva_dfm_1, sigmoid_table_71_0_sva_dfm_1,
          sigmoid_table_72_0_sva_dfm_1, sigmoid_table_73_0_sva_dfm_1, sigmoid_table_74_0_sva_dfm_1,
          sigmoid_table_75_0_sva_dfm_1, sigmoid_table_76_0_sva_dfm_1, sigmoid_table_77_0_sva_dfm_1,
          sigmoid_table_78_0_sva_dfm_1, sigmoid_table_79_0_sva_dfm_1, sigmoid_table_80_0_sva_dfm_1,
          sigmoid_table_81_0_sva_dfm_1, sigmoid_table_82_0_sva_dfm_1, sigmoid_table_83_0_sva_dfm_1,
          sigmoid_table_84_0_sva_dfm_1, sigmoid_table_85_0_sva_dfm_1, sigmoid_table_86_0_sva_dfm_1,
          sigmoid_table_87_0_sva_dfm_1, sigmoid_table_88_0_sva_dfm_1, sigmoid_table_89_0_sva_dfm_1,
          sigmoid_table_90_0_sva_dfm_1, sigmoid_table_91_0_sva_dfm_1, sigmoid_table_92_0_sva_dfm_1,
          sigmoid_table_93_0_sva_dfm_1, sigmoid_table_94_0_sva_dfm_1, sigmoid_table_95_0_sva_dfm_1,
          sigmoid_table_96_0_sva_dfm_1, sigmoid_table_97_0_sva_dfm_1, sigmoid_table_98_0_sva_dfm_1,
          sigmoid_table_99_0_sva_dfm_1, sigmoid_table_100_0_sva_dfm_1, sigmoid_table_101_0_sva_dfm_1,
          sigmoid_table_102_0_sva_dfm_1, sigmoid_table_103_0_sva_dfm_1, sigmoid_table_104_0_sva_dfm_1,
          sigmoid_table_105_0_sva_dfm_1, sigmoid_table_106_0_sva_dfm_1, sigmoid_table_107_0_sva_dfm_1,
          sigmoid_table_108_0_sva_dfm_1, sigmoid_table_109_0_sva_dfm_1, sigmoid_table_110_0_sva_dfm_1,
          sigmoid_table_111_0_sva_dfm_1, sigmoid_table_112_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          sigmoid_table_139_0_sva_dfm_1, sigmoid_table_140_0_sva_dfm_1, sigmoid_table_141_0_sva_dfm_1,
          sigmoid_table_142_0_sva_dfm_1, sigmoid_table_143_0_sva_dfm_1, sigmoid_table_144_0_sva_dfm_1,
          sigmoid_table_145_0_sva_dfm_1, sigmoid_table_146_0_sva_dfm_1, sigmoid_table_147_0_sva_dfm_1,
          sigmoid_table_148_0_sva_dfm_1, sigmoid_table_149_0_sva_dfm_1, sigmoid_table_150_0_sva_dfm_1,
          sigmoid_table_151_0_sva_dfm_1, sigmoid_table_152_0_sva_dfm_1, sigmoid_table_153_0_sva_dfm_1,
          sigmoid_table_154_0_sva_dfm_1, sigmoid_table_155_0_sva_dfm_1, sigmoid_table_156_0_sva_dfm_1,
          sigmoid_table_157_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_172_0_sva_dfm_1,
          sigmoid_table_173_0_sva_dfm_1, sigmoid_table_174_0_sva_dfm_1, sigmoid_table_175_0_sva_dfm_1,
          sigmoid_table_176_0_sva_dfm_1, sigmoid_table_177_0_sva_dfm_1, sigmoid_table_178_0_sva_dfm_1,
          sigmoid_table_179_0_sva_dfm_1, sigmoid_table_180_0_sva_dfm_1, sigmoid_table_181_0_sva_dfm_1,
          sigmoid_table_182_0_sva_dfm_1, sigmoid_table_183_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_194_0_sva_dfm_1,
          sigmoid_table_195_0_sva_dfm_1, sigmoid_table_196_0_sva_dfm_1, sigmoid_table_197_0_sva_dfm_1,
          sigmoid_table_198_0_sva_dfm_1, sigmoid_table_199_0_sva_dfm_1, sigmoid_table_200_0_sva_dfm_1,
          sigmoid_table_201_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, sigmoid_table_210_0_sva_dfm_1, sigmoid_table_211_0_sva_dfm_1, sigmoid_table_212_0_sva_dfm_1,
          sigmoid_table_213_0_sva_dfm_1, sigmoid_table_214_0_sva_dfm_1, sigmoid_table_215_0_sva_dfm_1,
          sigmoid_table_216_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_223_0_sva_dfm_1,
          sigmoid_table_224_0_sva_dfm_1, sigmoid_table_225_0_sva_dfm_1, sigmoid_table_226_0_sva_dfm_1,
          sigmoid_table_227_0_sva_dfm_1, sigmoid_table_228_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, sigmoid_table_234_0_sva_dfm_1, sigmoid_table_235_0_sva_dfm_1,
          sigmoid_table_236_0_sva_dfm_1, sigmoid_table_237_0_sva_dfm_1, sigmoid_table_238_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_243_0_sva_dfm_1, sigmoid_table_244_0_sva_dfm_1,
          sigmoid_table_245_0_sva_dfm_1, sigmoid_table_246_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_251_0_sva_dfm_1, sigmoid_table_252_0_sva_dfm_1,
          sigmoid_table_253_0_sva_dfm_1, sigmoid_table_254_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_259_0_sva_dfm_1, sigmoid_table_260_0_sva_dfm_1,
          sigmoid_table_261_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, sigmoid_table_265_0_sva_dfm_1,
          sigmoid_table_266_0_sva_dfm_1, sigmoid_table_267_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, sigmoid_table_271_0_sva_dfm_1, sigmoid_table_272_0_sva_dfm_1, sigmoid_table_273_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_276_0_sva_dfm_1, sigmoid_table_277_0_sva_dfm_1,
          sigmoid_table_278_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, sigmoid_table_282_0_sva_dfm_1,
          sigmoid_table_283_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_286_0_sva_dfm_1,
          sigmoid_table_287_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, sigmoid_table_291_0_sva_dfm_1,
          sigmoid_table_292_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_295_0_sva_dfm_1,
          sigmoid_table_296_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_299_0_sva_dfm_1,
          sigmoid_table_300_0_sva_dfm_1, 1'b0, sigmoid_table_302_0_sva_dfm_1, sigmoid_table_303_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_306_0_sva_dfm_1, sigmoid_table_307_0_sva_dfm_1,
          1'b0, sigmoid_table_309_0_sva_dfm_1, sigmoid_table_310_0_sva_dfm_1, 1'b0,
          sigmoid_table_312_0_sva_dfm_1, sigmoid_table_313_0_sva_dfm_1, 1'b0, sigmoid_table_315_0_sva_dfm_1,
          sigmoid_table_316_0_sva_dfm_1, 1'b0, sigmoid_table_318_0_sva_dfm_1, sigmoid_table_319_0_sva_dfm_1,
          1'b0, sigmoid_table_321_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_324_0_sva_dfm_1,
          1'b0, sigmoid_table_326_0_sva_dfm_1, sigmoid_table_327_0_sva_dfm_1, 1'b0,
          sigmoid_table_329_0_sva_dfm_1, 1'b0, sigmoid_table_331_0_sva_dfm_1, 1'b0,
          1'b0, sigmoid_table_334_0_sva_dfm_1, 1'b0, sigmoid_table_336_0_sva_dfm_1,
          1'b0, sigmoid_table_338_0_sva_dfm_1, 1'b0, sigmoid_table_340_0_sva_dfm_1,
          1'b0, sigmoid_table_342_0_sva_dfm_1, 1'b0, sigmoid_table_344_0_sva_dfm_1,
          1'b0, sigmoid_table_346_0_sva_dfm_1, 1'b0, sigmoid_table_348_0_sva_dfm_1,
          1'b0, sigmoid_table_350_0_sva_dfm_1, 1'b0, sigmoid_table_352_0_sva_dfm_1,
          1'b0, sigmoid_table_354_0_sva_dfm_1, sigmoid_table_355_0_sva_dfm_1, 1'b0,
          sigmoid_table_357_0_sva_dfm_1, 1'b0, sigmoid_table_359_0_sva_dfm_1, sigmoid_table_360_0_sva_dfm_1,
          1'b0, sigmoid_table_362_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_365_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_368_0_sva_dfm_1, sigmoid_table_369_0_sva_dfm_1,
          1'b0, sigmoid_table_371_0_sva_dfm_1, sigmoid_table_372_0_sva_dfm_1, 1'b0,
          1'b0, sigmoid_table_375_0_sva_dfm_1, sigmoid_table_376_0_sva_dfm_1, 1'b0,
          1'b0, sigmoid_table_379_0_sva_dfm_1, sigmoid_table_380_0_sva_dfm_1, sigmoid_table_381_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, sigmoid_table_385_0_sva_dfm_1, sigmoid_table_386_0_sva_dfm_1,
          sigmoid_table_387_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_394_0_sva_dfm_1,
          sigmoid_table_395_0_sva_dfm_1, sigmoid_table_396_0_sva_dfm_1, sigmoid_table_397_0_sva_dfm_1,
          sigmoid_table_398_0_sva_dfm_1, sigmoid_table_399_0_sva_dfm_1, sigmoid_table_400_0_sva_dfm_1,
          sigmoid_table_401_0_sva_dfm_1, sigmoid_table_402_0_sva_dfm_1, sigmoid_table_403_0_sva_dfm_1,
          sigmoid_table_404_0_sva_dfm_1, sigmoid_table_405_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, sigmoid_table_411_0_sva_dfm_1, sigmoid_table_412_0_sva_dfm_1,
          sigmoid_table_413_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, sigmoid_table_417_0_sva_dfm_1,
          sigmoid_table_418_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_421_0_sva_dfm_1,
          sigmoid_table_422_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_425_0_sva_dfm_1,
          sigmoid_table_426_0_sva_dfm_1, 1'b0, sigmoid_table_428_0_sva_dfm_1, sigmoid_table_429_0_sva_dfm_1,
          1'b0, sigmoid_table_431_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_434_0_sva_dfm_1,
          1'b0, sigmoid_table_436_0_sva_dfm_1, 1'b0, sigmoid_table_438_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_441_0_sva_dfm_1, 1'b0, sigmoid_table_443_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_446_0_sva_dfm_1, 1'b0, sigmoid_table_448_0_sva_dfm_1,
          1'b0, sigmoid_table_450_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_453_0_sva_dfm_1,
          1'b0, sigmoid_table_455_0_sva_dfm_1, sigmoid_table_456_0_sva_dfm_1, 1'b0,
          sigmoid_table_458_0_sva_dfm_1, sigmoid_table_459_0_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_462_0_sva_dfm_1, sigmoid_table_463_0_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_466_0_sva_dfm_1, sigmoid_table_467_0_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_470_0_sva_dfm_1, sigmoid_table_471_0_sva_dfm_1, sigmoid_table_472_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_475_0_sva_dfm_1, sigmoid_table_476_0_sva_dfm_1,
          sigmoid_table_477_0_sva_dfm_1, sigmoid_table_478_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_483_0_sva_dfm_1, sigmoid_table_484_0_sva_dfm_1,
          sigmoid_table_485_0_sva_dfm_1, sigmoid_table_486_0_sva_dfm_1, sigmoid_table_487_0_sva_dfm_1,
          sigmoid_table_488_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_516_0_sva_dfm_1,
          sigmoid_table_517_0_sva_dfm_1, sigmoid_table_518_0_sva_dfm_1, sigmoid_table_519_0_sva_dfm_1,
          sigmoid_table_520_0_sva_dfm_1, sigmoid_table_521_0_sva_dfm_1, sigmoid_table_522_0_sva_dfm_1,
          sigmoid_table_523_0_sva_dfm_1, sigmoid_table_524_0_sva_dfm_1, sigmoid_table_525_0_sva_dfm_1,
          sigmoid_table_526_0_sva_dfm_1, sigmoid_table_527_0_sva_dfm_1, sigmoid_table_528_0_sva_dfm_1,
          sigmoid_table_529_0_sva_dfm_1, sigmoid_table_530_0_sva_dfm_1, sigmoid_table_531_0_sva_dfm_1,
          sigmoid_table_532_0_sva_dfm_1, sigmoid_table_533_0_sva_dfm_1, sigmoid_table_534_0_sva_dfm_1,
          sigmoid_table_535_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_542_0_sva_dfm_1,
          sigmoid_table_543_0_sva_dfm_1, sigmoid_table_544_0_sva_dfm_1, sigmoid_table_545_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_550_0_sva_dfm_1, sigmoid_table_551_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, sigmoid_table_555_0_sva_dfm_1, sigmoid_table_556_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_559_0_sva_dfm_1, sigmoid_table_560_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_563_0_sva_dfm_1, sigmoid_table_564_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_567_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_570_0_sva_dfm_1,
          1'b0, sigmoid_table_572_0_sva_dfm_1, sigmoid_table_573_0_sva_dfm_1, 1'b0,
          sigmoid_table_575_0_sva_dfm_1, 1'b0, sigmoid_table_577_0_sva_dfm_1, 1'b0,
          sigmoid_table_579_0_sva_dfm_1, sigmoid_table_580_0_sva_dfm_1, 1'b0, sigmoid_table_582_0_sva_dfm_1,
          1'b0, sigmoid_table_584_0_sva_dfm_1, sigmoid_table_585_0_sva_dfm_1, 1'b0,
          sigmoid_table_587_0_sva_dfm_1, 1'b0, sigmoid_table_589_0_sva_dfm_1, 1'b0,
          sigmoid_table_591_0_sva_dfm_1, sigmoid_table_592_0_sva_dfm_1, 1'b0, sigmoid_table_594_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_597_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_600_0_sva_dfm_1,
          sigmoid_table_601_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_604_0_sva_dfm_1,
          sigmoid_table_605_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_608_0_sva_dfm_1,
          sigmoid_table_609_0_sva_dfm_1, sigmoid_table_610_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, sigmoid_table_614_0_sva_dfm_1, sigmoid_table_615_0_sva_dfm_1, sigmoid_table_616_0_sva_dfm_1,
          sigmoid_table_617_0_sva_dfm_1, sigmoid_table_618_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_631_0_sva_dfm_1,
          sigmoid_table_632_0_sva_dfm_1, sigmoid_table_633_0_sva_dfm_1, sigmoid_table_634_0_sva_dfm_1,
          sigmoid_table_635_0_sva_dfm_1, sigmoid_table_636_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, sigmoid_table_640_0_sva_dfm_1, sigmoid_table_641_0_sva_dfm_1, sigmoid_table_642_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, sigmoid_table_646_0_sva_dfm_1, sigmoid_table_647_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_650_0_sva_dfm_1, sigmoid_table_651_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_654_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_657_0_sva_dfm_1,
          sigmoid_table_658_0_sva_dfm_1, 1'b0, sigmoid_table_660_0_sva_dfm_1, sigmoid_table_661_0_sva_dfm_1,
          1'b0, sigmoid_table_663_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_666_0_sva_dfm_1,
          1'b0, sigmoid_table_668_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_671_0_sva_dfm_1,
          1'b0, sigmoid_table_673_0_sva_dfm_1, 1'b0, sigmoid_table_675_0_sva_dfm_1,
          1'b0, sigmoid_table_677_0_sva_dfm_1, 1'b0, sigmoid_table_679_0_sva_dfm_1,
          1'b0, sigmoid_table_681_0_sva_dfm_1, 1'b0, sigmoid_table_683_0_sva_dfm_1,
          1'b0, sigmoid_table_685_0_sva_dfm_1, 1'b0, sigmoid_table_687_0_sva_dfm_1,
          1'b0, sigmoid_table_689_0_sva_dfm_1, 1'b0, sigmoid_table_691_0_sva_dfm_1,
          sigmoid_table_692_0_sva_dfm_1, 1'b0, sigmoid_table_694_0_sva_dfm_1, 1'b0,
          sigmoid_table_696_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_699_0_sva_dfm_1,
          1'b0, sigmoid_table_701_0_sva_dfm_1, sigmoid_table_702_0_sva_dfm_1, 1'b0,
          sigmoid_table_704_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_707_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_710_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_713_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_716_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_719_0_sva_dfm_1,
          sigmoid_table_720_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_723_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_726_0_sva_dfm_1, sigmoid_table_727_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_730_0_sva_dfm_1, sigmoid_table_731_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_734_0_sva_dfm_1, sigmoid_table_735_0_sva_dfm_1,
          sigmoid_table_736_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_739_0_sva_dfm_1,
          sigmoid_table_740_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_743_0_sva_dfm_1,
          sigmoid_table_744_0_sva_dfm_1, sigmoid_table_745_0_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_748_0_sva_dfm_1, sigmoid_table_749_0_sva_dfm_1, sigmoid_table_750_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, sigmoid_table_754_0_sva_dfm_1, sigmoid_table_755_0_sva_dfm_1,
          sigmoid_table_756_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, sigmoid_table_760_0_sva_dfm_1,
          sigmoid_table_761_0_sva_dfm_1, sigmoid_table_762_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, sigmoid_table_766_0_sva_dfm_1, sigmoid_table_767_0_sva_dfm_1, sigmoid_table_768_0_sva_dfm_1,
          sigmoid_table_769_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_774_0_sva_dfm_1,
          sigmoid_table_775_0_sva_dfm_1, sigmoid_table_776_0_sva_dfm_1, sigmoid_table_777_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_782_0_sva_dfm_1, sigmoid_table_783_0_sva_dfm_1,
          sigmoid_table_784_0_sva_dfm_1, sigmoid_table_785_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, sigmoid_table_791_0_sva_dfm_1, sigmoid_table_792_0_sva_dfm_1,
          sigmoid_table_793_0_sva_dfm_1, sigmoid_table_794_0_sva_dfm_1, sigmoid_table_795_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_802_0_sva_dfm_1, sigmoid_table_803_0_sva_dfm_1,
          sigmoid_table_804_0_sva_dfm_1, sigmoid_table_805_0_sva_dfm_1, sigmoid_table_806_0_sva_dfm_1,
          sigmoid_table_807_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          sigmoid_table_815_0_sva_dfm_1, sigmoid_table_816_0_sva_dfm_1, sigmoid_table_817_0_sva_dfm_1,
          sigmoid_table_818_0_sva_dfm_1, sigmoid_table_819_0_sva_dfm_1, sigmoid_table_820_0_sva_dfm_1,
          sigmoid_table_821_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_831_0_sva_dfm_1, sigmoid_table_832_0_sva_dfm_1,
          sigmoid_table_833_0_sva_dfm_1, sigmoid_table_834_0_sva_dfm_1, sigmoid_table_835_0_sva_dfm_1,
          sigmoid_table_836_0_sva_dfm_1, sigmoid_table_837_0_sva_dfm_1, sigmoid_table_838_0_sva_dfm_1,
          sigmoid_table_839_0_sva_dfm_1, sigmoid_table_840_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_853_0_sva_dfm_1,
          sigmoid_table_854_0_sva_dfm_1, sigmoid_table_855_0_sva_dfm_1, sigmoid_table_856_0_sva_dfm_1,
          sigmoid_table_857_0_sva_dfm_1, sigmoid_table_858_0_sva_dfm_1, sigmoid_table_859_0_sva_dfm_1,
          sigmoid_table_860_0_sva_dfm_1, sigmoid_table_861_0_sva_dfm_1, sigmoid_table_862_0_sva_dfm_1,
          sigmoid_table_863_0_sva_dfm_1, sigmoid_table_864_0_sva_dfm_1, sigmoid_table_865_0_sva_dfm_1,
          sigmoid_table_866_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_885_0_sva_dfm_1,
          sigmoid_table_886_0_sva_dfm_1, sigmoid_table_887_0_sva_dfm_1, sigmoid_table_888_0_sva_dfm_1,
          sigmoid_table_889_0_sva_dfm_1, sigmoid_table_890_0_sva_dfm_1, sigmoid_table_891_0_sva_dfm_1,
          sigmoid_table_892_0_sva_dfm_1, sigmoid_table_893_0_sva_dfm_1, sigmoid_table_894_0_sva_dfm_1,
          sigmoid_table_895_0_sva_dfm_1, sigmoid_table_896_0_sva_dfm_1, sigmoid_table_897_0_sva_dfm_1,
          sigmoid_table_898_0_sva_dfm_1, sigmoid_table_899_0_sva_dfm_1, sigmoid_table_900_0_sva_dfm_1,
          sigmoid_table_901_0_sva_dfm_1, sigmoid_table_902_0_sva_dfm_1, sigmoid_table_903_0_sva_dfm_1,
          sigmoid_table_904_0_sva_dfm_1, sigmoid_table_905_0_sva_dfm_1, sigmoid_table_906_0_sva_dfm_1,
          sigmoid_table_907_0_sva_dfm_1, sigmoid_table_908_0_sva_dfm_1, sigmoid_table_909_0_sva_dfm_1,
          sigmoid_table_910_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, sigmoid_table_955_0_sva_dfm_1, sigmoid_table_956_0_sva_dfm_1, sigmoid_table_957_0_sva_dfm_1,
          sigmoid_table_958_0_sva_dfm_1, sigmoid_table_959_0_sva_dfm_1, sigmoid_table_960_0_sva_dfm_1,
          sigmoid_table_961_0_sva_dfm_1, sigmoid_table_962_0_sva_dfm_1, sigmoid_table_963_0_sva_dfm_1,
          sigmoid_table_964_0_sva_dfm_1, sigmoid_table_965_0_sva_dfm_1, sigmoid_table_966_0_sva_dfm_1,
          sigmoid_table_967_0_sva_dfm_1, sigmoid_table_968_0_sva_dfm_1, sigmoid_table_969_0_sva_dfm_1,
          sigmoid_table_970_0_sva_dfm_1, sigmoid_table_971_0_sva_dfm_1, sigmoid_table_972_0_sva_dfm_1,
          sigmoid_table_973_0_sva_dfm_1, sigmoid_table_974_0_sva_dfm_1, sigmoid_table_975_0_sva_dfm_1,
          sigmoid_table_976_0_sva_dfm_1, sigmoid_table_977_0_sva_dfm_1, sigmoid_table_978_0_sva_dfm_1,
          sigmoid_table_979_0_sva_dfm_1, sigmoid_table_980_0_sva_dfm_1, sigmoid_table_981_0_sva_dfm_1,
          sigmoid_table_982_0_sva_dfm_1, sigmoid_table_983_0_sva_dfm_1, sigmoid_table_984_0_sva_dfm_1,
          sigmoid_table_985_0_sva_dfm_1, sigmoid_table_986_0_sva_dfm_1, sigmoid_table_987_0_sva_dfm_1,
          sigmoid_table_988_0_sva_dfm_1, sigmoid_table_989_0_sva_dfm_1, sigmoid_table_990_0_sva_dfm_1,
          sigmoid_table_991_0_sva_dfm_1, sigmoid_table_992_0_sva_dfm_1, sigmoid_table_993_0_sva_dfm_1,
          sigmoid_table_994_0_sva_dfm_1, sigmoid_table_995_0_sva_dfm_1, sigmoid_table_996_0_sva_dfm_1,
          sigmoid_table_997_0_sva_dfm_1, sigmoid_table_998_0_sva_dfm_1, sigmoid_table_999_0_sva_dfm_1,
          sigmoid_table_1000_0_sva_dfm_1, sigmoid_table_1001_0_sva_dfm_1, sigmoid_table_1002_0_sva_dfm_1,
          sigmoid_table_1003_0_sva_dfm_1, sigmoid_table_1004_0_sva_dfm_1, sigmoid_table_1005_0_sva_dfm_1,
          sigmoid_table_1006_0_sva_dfm_1, sigmoid_table_1007_0_sva_dfm_1, sigmoid_table_1008_0_sva_dfm_1,
          sigmoid_table_1009_0_sva_dfm_1, sigmoid_table_1010_0_sva_dfm_1, sigmoid_table_1011_0_sva_dfm_1,
          sigmoid_table_1012_0_sva_dfm_1, sigmoid_table_1013_0_sva_dfm_1, sigmoid_table_1014_0_sva_dfm_1,
          sigmoid_table_1015_0_sva_dfm_1, sigmoid_table_1016_0_sva_dfm_1, sigmoid_table_1017_0_sva_dfm_1,
          sigmoid_table_1018_0_sva_dfm_1, sigmoid_table_1019_0_sva_dfm_1, sigmoid_table_1020_0_sva_dfm_1,
          sigmoid_table_1021_0_sva_dfm_1, sigmoid_table_1022_0_sva_dfm_1, sigmoid_table_1023_0_sva_dfm_1,
          {for_for_or_1_itm , for_for_or_itm});
      res_rsci_d_9 <= MUX_s_1_1024_2(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          sigmoid_table_512_9_sva_dfm_1, sigmoid_table_513_9_sva_dfm_1, sigmoid_table_514_9_sva_dfm_1,
          sigmoid_table_515_9_sva_dfm_1, sigmoid_table_516_9_sva_dfm_1, sigmoid_table_517_9_sva_dfm_1,
          sigmoid_table_518_9_sva_dfm_1, sigmoid_table_519_9_sva_dfm_1, sigmoid_table_520_9_sva_dfm_1,
          sigmoid_table_521_9_sva_dfm_1, sigmoid_table_522_9_sva_dfm_1, sigmoid_table_523_9_sva_dfm_1,
          sigmoid_table_524_9_sva_dfm_1, sigmoid_table_525_9_sva_dfm_1, sigmoid_table_526_9_sva_dfm_1,
          sigmoid_table_527_9_sva_dfm_1, sigmoid_table_528_9_sva_dfm_1, sigmoid_table_529_9_sva_dfm_1,
          sigmoid_table_530_9_sva_dfm_1, sigmoid_table_531_9_sva_dfm_1, sigmoid_table_532_9_sva_dfm_1,
          sigmoid_table_533_9_sva_dfm_1, sigmoid_table_534_9_sva_dfm_1, sigmoid_table_535_9_sva_dfm_1,
          sigmoid_table_536_9_sva_dfm_1, sigmoid_table_537_9_sva_dfm_1, sigmoid_table_538_9_sva_dfm_1,
          sigmoid_table_539_9_sva_dfm_1, sigmoid_table_540_9_sva_dfm_1, sigmoid_table_541_9_sva_dfm_1,
          sigmoid_table_542_9_sva_dfm_1, sigmoid_table_543_9_sva_dfm_1, sigmoid_table_544_9_sva_dfm_1,
          sigmoid_table_545_9_sva_dfm_1, sigmoid_table_546_9_sva_dfm_1, sigmoid_table_547_9_sva_dfm_1,
          sigmoid_table_548_9_sva_dfm_1, sigmoid_table_549_9_sva_dfm_1, sigmoid_table_550_9_sva_dfm_1,
          sigmoid_table_551_9_sva_dfm_1, sigmoid_table_552_9_sva_dfm_1, sigmoid_table_553_9_sva_dfm_1,
          sigmoid_table_554_9_sva_dfm_1, sigmoid_table_555_9_sva_dfm_1, sigmoid_table_556_9_sva_dfm_1,
          sigmoid_table_557_9_sva_dfm_1, sigmoid_table_558_9_sva_dfm_1, sigmoid_table_559_9_sva_dfm_1,
          sigmoid_table_560_9_sva_dfm_1, sigmoid_table_561_9_sva_dfm_1, sigmoid_table_562_9_sva_dfm_1,
          sigmoid_table_563_9_sva_dfm_1, sigmoid_table_564_9_sva_dfm_1, sigmoid_table_565_9_sva_dfm_1,
          sigmoid_table_566_9_sva_dfm_1, sigmoid_table_567_9_sva_dfm_1, sigmoid_table_568_9_sva_dfm_1,
          sigmoid_table_569_9_sva_dfm_1, sigmoid_table_570_9_sva_dfm_1, sigmoid_table_571_9_sva_dfm_1,
          sigmoid_table_572_9_sva_dfm_1, sigmoid_table_573_9_sva_dfm_1, sigmoid_table_574_9_sva_dfm_1,
          sigmoid_table_575_9_sva_dfm_1, sigmoid_table_576_9_sva_dfm_1, sigmoid_table_577_9_sva_dfm_1,
          sigmoid_table_578_9_sva_dfm_1, sigmoid_table_579_9_sva_dfm_1, sigmoid_table_580_9_sva_dfm_1,
          sigmoid_table_581_9_sva_dfm_1, sigmoid_table_582_9_sva_dfm_1, sigmoid_table_583_8_sva_dfm_1,
          sigmoid_table_584_8_sva_dfm_1, sigmoid_table_585_8_sva_dfm_1, sigmoid_table_586_8_sva_dfm_1,
          sigmoid_table_587_8_sva_dfm_1, sigmoid_table_588_8_sva_dfm_1, sigmoid_table_589_8_sva_dfm_1,
          sigmoid_table_590_8_sva_dfm_1, sigmoid_table_591_8_sva_dfm_1, sigmoid_table_592_8_sva_dfm_1,
          sigmoid_table_593_8_sva_dfm_1, sigmoid_table_594_8_sva_dfm_1, sigmoid_table_595_8_sva_dfm_1,
          sigmoid_table_596_8_sva_dfm_1, sigmoid_table_597_8_sva_dfm_1, sigmoid_table_598_8_sva_dfm_1,
          sigmoid_table_599_8_sva_dfm_1, sigmoid_table_600_8_sva_dfm_1, sigmoid_table_601_8_sva_dfm_1,
          sigmoid_table_602_8_sva_dfm_1, sigmoid_table_603_8_sva_dfm_1, sigmoid_table_604_8_sva_dfm_1,
          sigmoid_table_605_8_sva_dfm_1, sigmoid_table_606_8_sva_dfm_1, sigmoid_table_607_8_sva_dfm_1,
          sigmoid_table_608_8_sva_dfm_1, sigmoid_table_609_8_sva_dfm_1, sigmoid_table_610_8_sva_dfm_1,
          sigmoid_table_611_8_sva_dfm_1, sigmoid_table_612_8_sva_dfm_1, sigmoid_table_613_8_sva_dfm_1,
          sigmoid_table_614_8_sva_dfm_1, sigmoid_table_615_8_sva_dfm_1, sigmoid_table_616_8_sva_dfm_1,
          sigmoid_table_617_8_sva_dfm_1, sigmoid_table_618_8_sva_dfm_1, sigmoid_table_619_8_sva_dfm_1,
          sigmoid_table_620_8_sva_dfm_1, sigmoid_table_621_8_sva_dfm_1, sigmoid_table_622_8_sva_dfm_1,
          sigmoid_table_623_8_sva_dfm_1, sigmoid_table_624_8_sva_dfm_1, sigmoid_table_625_8_sva_dfm_1,
          sigmoid_table_626_8_sva_dfm_1, sigmoid_table_627_8_sva_dfm_1, sigmoid_table_628_8_sva_dfm_1,
          sigmoid_table_629_8_sva_dfm_1, sigmoid_table_630_8_sva_dfm_1, sigmoid_table_631_8_sva_dfm_1,
          sigmoid_table_632_8_sva_dfm_1, sigmoid_table_633_8_sva_dfm_1, sigmoid_table_634_8_sva_dfm_1,
          sigmoid_table_635_8_sva_dfm_1, sigmoid_table_636_8_sva_dfm_1, sigmoid_table_637_7_sva_dfm_1,
          sigmoid_table_638_7_sva_dfm_1, sigmoid_table_639_7_sva_dfm_1, sigmoid_table_640_7_sva_dfm_1,
          sigmoid_table_641_7_sva_dfm_1, sigmoid_table_642_7_sva_dfm_1, sigmoid_table_643_7_sva_dfm_1,
          sigmoid_table_644_7_sva_dfm_1, sigmoid_table_645_7_sva_dfm_1, sigmoid_table_646_7_sva_dfm_1,
          sigmoid_table_647_7_sva_dfm_1, sigmoid_table_648_7_sva_dfm_1, sigmoid_table_649_7_sva_dfm_1,
          sigmoid_table_650_7_sva_dfm_1, sigmoid_table_651_7_sva_dfm_1, sigmoid_table_652_7_sva_dfm_1,
          sigmoid_table_653_7_sva_dfm_1, sigmoid_table_654_7_sva_dfm_1, sigmoid_table_655_7_sva_dfm_1,
          sigmoid_table_656_7_sva_dfm_1, sigmoid_table_657_7_sva_dfm_1, sigmoid_table_658_7_sva_dfm_1,
          sigmoid_table_659_7_sva_dfm_1, sigmoid_table_660_7_sva_dfm_1, sigmoid_table_661_7_sva_dfm_1,
          sigmoid_table_662_7_sva_dfm_1, sigmoid_table_663_7_sva_dfm_1, sigmoid_table_664_7_sva_dfm_1,
          sigmoid_table_665_7_sva_dfm_1, sigmoid_table_666_7_sva_dfm_1, sigmoid_table_667_7_sva_dfm_1,
          sigmoid_table_668_7_sva_dfm_1, sigmoid_table_669_7_sva_dfm_1, sigmoid_table_670_7_sva_dfm_1,
          sigmoid_table_671_7_sva_dfm_1, sigmoid_table_672_7_sva_dfm_1, sigmoid_table_673_7_sva_dfm_1,
          sigmoid_table_674_7_sva_dfm_1, sigmoid_table_675_7_sva_dfm_1, sigmoid_table_676_7_sva_dfm_1,
          sigmoid_table_677_7_sva_dfm_1, sigmoid_table_678_7_sva_dfm_1, sigmoid_table_679_7_sva_dfm_1,
          sigmoid_table_680_7_sva_dfm_1, sigmoid_table_681_7_sva_dfm_1, sigmoid_table_682_7_sva_dfm_1,
          sigmoid_table_683_7_sva_dfm_1, sigmoid_table_684_7_sva_dfm_1, sigmoid_table_685_7_sva_dfm_1,
          sigmoid_table_686_6_sva_dfm_1, sigmoid_table_687_6_sva_dfm_1, sigmoid_table_688_6_sva_dfm_1,
          sigmoid_table_689_6_sva_dfm_1, sigmoid_table_690_6_sva_dfm_1, sigmoid_table_691_6_sva_dfm_1,
          sigmoid_table_692_6_sva_dfm_1, sigmoid_table_693_6_sva_dfm_1, sigmoid_table_694_6_sva_dfm_1,
          sigmoid_table_695_6_sva_dfm_1, sigmoid_table_696_6_sva_dfm_1, sigmoid_table_697_6_sva_dfm_1,
          sigmoid_table_698_6_sva_dfm_1, sigmoid_table_699_6_sva_dfm_1, sigmoid_table_700_6_sva_dfm_1,
          sigmoid_table_701_6_sva_dfm_1, sigmoid_table_702_6_sva_dfm_1, sigmoid_table_703_6_sva_dfm_1,
          sigmoid_table_704_6_sva_dfm_1, sigmoid_table_705_6_sva_dfm_1, sigmoid_table_706_6_sva_dfm_1,
          sigmoid_table_707_6_sva_dfm_1, sigmoid_table_708_6_sva_dfm_1, sigmoid_table_709_6_sva_dfm_1,
          sigmoid_table_710_6_sva_dfm_1, sigmoid_table_711_6_sva_dfm_1, sigmoid_table_712_6_sva_dfm_1,
          sigmoid_table_713_6_sva_dfm_1, sigmoid_table_714_6_sva_dfm_1, sigmoid_table_715_6_sva_dfm_1,
          sigmoid_table_716_6_sva_dfm_1, sigmoid_table_717_6_sva_dfm_1, sigmoid_table_718_6_sva_dfm_1,
          sigmoid_table_719_6_sva_dfm_1, sigmoid_table_720_6_sva_dfm_1, sigmoid_table_721_6_sva_dfm_1,
          sigmoid_table_722_6_sva_dfm_1, sigmoid_table_723_6_sva_dfm_1, sigmoid_table_724_6_sva_dfm_1,
          sigmoid_table_725_6_sva_dfm_1, sigmoid_table_726_6_sva_dfm_1, sigmoid_table_727_6_sva_dfm_1,
          sigmoid_table_728_6_sva_dfm_1, sigmoid_table_729_6_sva_dfm_1, sigmoid_table_730_6_sva_dfm_1,
          sigmoid_table_731_6_sva_dfm_1, sigmoid_table_732_5_sva_dfm_1, sigmoid_table_733_5_sva_dfm_1,
          sigmoid_table_734_5_sva_dfm_1, sigmoid_table_735_5_sva_dfm_1, sigmoid_table_736_5_sva_dfm_1,
          sigmoid_table_737_5_sva_dfm_1, sigmoid_table_738_5_sva_dfm_1, sigmoid_table_739_5_sva_dfm_1,
          sigmoid_table_740_5_sva_dfm_1, sigmoid_table_741_5_sva_dfm_1, sigmoid_table_742_5_sva_dfm_1,
          sigmoid_table_743_5_sva_dfm_1, sigmoid_table_744_5_sva_dfm_1, sigmoid_table_745_5_sva_dfm_1,
          sigmoid_table_746_5_sva_dfm_1, sigmoid_table_747_5_sva_dfm_1, sigmoid_table_748_5_sva_dfm_1,
          sigmoid_table_749_5_sva_dfm_1, sigmoid_table_750_5_sva_dfm_1, sigmoid_table_751_5_sva_dfm_1,
          sigmoid_table_752_5_sva_dfm_1, sigmoid_table_753_5_sva_dfm_1, sigmoid_table_754_5_sva_dfm_1,
          sigmoid_table_755_5_sva_dfm_1, sigmoid_table_756_5_sva_dfm_1, sigmoid_table_757_5_sva_dfm_1,
          sigmoid_table_758_5_sva_dfm_1, sigmoid_table_759_5_sva_dfm_1, sigmoid_table_760_5_sva_dfm_1,
          sigmoid_table_761_5_sva_dfm_1, sigmoid_table_762_5_sva_dfm_1, sigmoid_table_763_5_sva_dfm_1,
          sigmoid_table_764_5_sva_dfm_1, sigmoid_table_765_5_sva_dfm_1, sigmoid_table_766_5_sva_dfm_1,
          sigmoid_table_767_5_sva_dfm_1, sigmoid_table_768_5_sva_dfm_1, sigmoid_table_769_5_sva_dfm_1,
          sigmoid_table_770_5_sva_dfm_1, sigmoid_table_771_5_sva_dfm_1, sigmoid_table_772_5_sva_dfm_1,
          sigmoid_table_773_5_sva_dfm_1, sigmoid_table_774_5_sva_dfm_1, sigmoid_table_775_5_sva_dfm_1,
          sigmoid_table_776_5_sva_dfm_1, sigmoid_table_777_5_sva_dfm_1, sigmoid_table_778_4_sva_dfm_1,
          sigmoid_table_779_4_sva_dfm_1, sigmoid_table_780_4_sva_dfm_1, sigmoid_table_781_4_sva_dfm_1,
          sigmoid_table_782_4_sva_dfm_1, sigmoid_table_783_4_sva_dfm_1, sigmoid_table_784_4_sva_dfm_1,
          sigmoid_table_785_4_sva_dfm_1, sigmoid_table_786_4_sva_dfm_1, sigmoid_table_787_4_sva_dfm_1,
          sigmoid_table_788_4_sva_dfm_1, sigmoid_table_789_4_sva_dfm_1, sigmoid_table_790_4_sva_dfm_1,
          sigmoid_table_791_4_sva_dfm_1, sigmoid_table_792_4_sva_dfm_1, sigmoid_table_793_4_sva_dfm_1,
          sigmoid_table_794_4_sva_dfm_1, sigmoid_table_795_4_sva_dfm_1, sigmoid_table_796_4_sva_dfm_1,
          sigmoid_table_797_4_sva_dfm_1, sigmoid_table_798_4_sva_dfm_1, sigmoid_table_799_4_sva_dfm_1,
          sigmoid_table_800_4_sva_dfm_1, sigmoid_table_801_4_sva_dfm_1, sigmoid_table_802_4_sva_dfm_1,
          sigmoid_table_803_4_sva_dfm_1, sigmoid_table_804_4_sva_dfm_1, sigmoid_table_805_4_sva_dfm_1,
          sigmoid_table_806_4_sva_dfm_1, sigmoid_table_807_4_sva_dfm_1, sigmoid_table_808_4_sva_dfm_1,
          sigmoid_table_809_4_sva_dfm_1, sigmoid_table_810_4_sva_dfm_1, sigmoid_table_811_4_sva_dfm_1,
          sigmoid_table_812_4_sva_dfm_1, sigmoid_table_813_4_sva_dfm_1, sigmoid_table_814_4_sva_dfm_1,
          sigmoid_table_815_4_sva_dfm_1, sigmoid_table_816_4_sva_dfm_1, sigmoid_table_817_4_sva_dfm_1,
          sigmoid_table_818_4_sva_dfm_1, sigmoid_table_819_4_sva_dfm_1, sigmoid_table_820_4_sva_dfm_1,
          sigmoid_table_821_4_sva_dfm_1, sigmoid_table_822_3_sva_dfm_1, sigmoid_table_823_3_sva_dfm_1,
          sigmoid_table_824_3_sva_dfm_1, sigmoid_table_825_3_sva_dfm_1, sigmoid_table_826_3_sva_dfm_1,
          sigmoid_table_827_3_sva_dfm_1, sigmoid_table_828_3_sva_dfm_1, sigmoid_table_829_3_sva_dfm_1,
          sigmoid_table_830_3_sva_dfm_1, sigmoid_table_831_3_sva_dfm_1, sigmoid_table_832_3_sva_dfm_1,
          sigmoid_table_833_3_sva_dfm_1, sigmoid_table_834_3_sva_dfm_1, sigmoid_table_835_3_sva_dfm_1,
          sigmoid_table_836_3_sva_dfm_1, sigmoid_table_837_3_sva_dfm_1, sigmoid_table_838_3_sva_dfm_1,
          sigmoid_table_839_3_sva_dfm_1, sigmoid_table_840_3_sva_dfm_1, sigmoid_table_841_3_sva_dfm_1,
          sigmoid_table_842_3_sva_dfm_1, sigmoid_table_843_3_sva_dfm_1, sigmoid_table_844_3_sva_dfm_1,
          sigmoid_table_845_3_sva_dfm_1, sigmoid_table_846_3_sva_dfm_1, sigmoid_table_847_3_sva_dfm_1,
          sigmoid_table_848_3_sva_dfm_1, sigmoid_table_849_3_sva_dfm_1, sigmoid_table_850_3_sva_dfm_1,
          sigmoid_table_851_3_sva_dfm_1, sigmoid_table_852_3_sva_dfm_1, sigmoid_table_853_3_sva_dfm_1,
          sigmoid_table_854_3_sva_dfm_1, sigmoid_table_855_3_sva_dfm_1, sigmoid_table_856_3_sva_dfm_1,
          sigmoid_table_857_3_sva_dfm_1, sigmoid_table_858_3_sva_dfm_1, sigmoid_table_859_3_sva_dfm_1,
          sigmoid_table_860_3_sva_dfm_1, sigmoid_table_861_3_sva_dfm_1, sigmoid_table_862_3_sva_dfm_1,
          sigmoid_table_863_3_sva_dfm_1, sigmoid_table_864_3_sva_dfm_1, sigmoid_table_865_3_sva_dfm_1,
          sigmoid_table_866_3_sva_dfm_1, sigmoid_table_867_2_sva_dfm_1, sigmoid_table_868_2_sva_dfm_1,
          sigmoid_table_869_2_sva_dfm_1, sigmoid_table_870_2_sva_dfm_1, sigmoid_table_871_2_sva_dfm_1,
          sigmoid_table_872_2_sva_dfm_1, sigmoid_table_873_2_sva_dfm_1, sigmoid_table_874_2_sva_dfm_1,
          sigmoid_table_875_2_sva_dfm_1, sigmoid_table_876_2_sva_dfm_1, sigmoid_table_877_2_sva_dfm_1,
          sigmoid_table_878_2_sva_dfm_1, sigmoid_table_879_2_sva_dfm_1, sigmoid_table_880_2_sva_dfm_1,
          sigmoid_table_881_2_sva_dfm_1, sigmoid_table_882_2_sva_dfm_1, sigmoid_table_883_2_sva_dfm_1,
          sigmoid_table_884_2_sva_dfm_1, sigmoid_table_885_2_sva_dfm_1, sigmoid_table_886_2_sva_dfm_1,
          sigmoid_table_887_2_sva_dfm_1, sigmoid_table_888_2_sva_dfm_1, sigmoid_table_889_2_sva_dfm_1,
          sigmoid_table_890_2_sva_dfm_1, sigmoid_table_891_2_sva_dfm_1, sigmoid_table_892_2_sva_dfm_1,
          sigmoid_table_893_2_sva_dfm_1, sigmoid_table_894_2_sva_dfm_1, sigmoid_table_895_2_sva_dfm_1,
          sigmoid_table_896_2_sva_dfm_1, sigmoid_table_897_2_sva_dfm_1, sigmoid_table_898_2_sva_dfm_1,
          sigmoid_table_899_2_sva_dfm_1, sigmoid_table_900_2_sva_dfm_1, sigmoid_table_901_2_sva_dfm_1,
          sigmoid_table_902_2_sva_dfm_1, sigmoid_table_903_2_sva_dfm_1, sigmoid_table_904_2_sva_dfm_1,
          sigmoid_table_905_2_sva_dfm_1, sigmoid_table_906_2_sva_dfm_1, sigmoid_table_907_2_sva_dfm_1,
          sigmoid_table_908_2_sva_dfm_1, sigmoid_table_909_2_sva_dfm_1, sigmoid_table_910_2_sva_dfm_1,
          sigmoid_table_911_1_sva_dfm_1, sigmoid_table_912_1_sva_dfm_1, sigmoid_table_913_1_sva_dfm_1,
          sigmoid_table_914_1_sva_dfm_1, sigmoid_table_915_1_sva_dfm_1, sigmoid_table_916_1_sva_dfm_1,
          sigmoid_table_917_1_sva_dfm_1, sigmoid_table_918_1_sva_dfm_1, sigmoid_table_919_1_sva_dfm_1,
          sigmoid_table_920_1_sva_dfm_1, sigmoid_table_921_1_sva_dfm_1, sigmoid_table_922_1_sva_dfm_1,
          sigmoid_table_923_1_sva_dfm_1, sigmoid_table_924_1_sva_dfm_1, sigmoid_table_925_1_sva_dfm_1,
          sigmoid_table_926_1_sva_dfm_1, sigmoid_table_927_1_sva_dfm_1, sigmoid_table_928_1_sva_dfm_1,
          sigmoid_table_929_1_sva_dfm_1, sigmoid_table_930_1_sva_dfm_1, sigmoid_table_931_1_sva_dfm_1,
          sigmoid_table_932_1_sva_dfm_1, sigmoid_table_933_1_sva_dfm_1, sigmoid_table_934_1_sva_dfm_1,
          sigmoid_table_935_1_sva_dfm_1, sigmoid_table_936_1_sva_dfm_1, sigmoid_table_937_1_sva_dfm_1,
          sigmoid_table_938_1_sva_dfm_1, sigmoid_table_939_1_sva_dfm_1, sigmoid_table_940_1_sva_dfm_1,
          sigmoid_table_941_1_sva_dfm_1, sigmoid_table_942_1_sva_dfm_1, sigmoid_table_943_1_sva_dfm_1,
          sigmoid_table_944_1_sva_dfm_1, sigmoid_table_945_1_sva_dfm_1, sigmoid_table_946_1_sva_dfm_1,
          sigmoid_table_947_1_sva_dfm_1, sigmoid_table_948_1_sva_dfm_1, sigmoid_table_949_1_sva_dfm_1,
          sigmoid_table_950_1_sva_dfm_1, sigmoid_table_951_1_sva_dfm_1, sigmoid_table_952_1_sva_dfm_1,
          sigmoid_table_953_1_sva_dfm_1, sigmoid_table_954_1_sva_dfm_1, sigmoid_table_955_0_sva_dfm_1,
          sigmoid_table_956_0_sva_dfm_1, sigmoid_table_957_0_sva_dfm_1, sigmoid_table_958_0_sva_dfm_1,
          sigmoid_table_959_0_sva_dfm_1, sigmoid_table_960_0_sva_dfm_1, sigmoid_table_961_0_sva_dfm_1,
          sigmoid_table_962_0_sva_dfm_1, sigmoid_table_963_0_sva_dfm_1, sigmoid_table_964_0_sva_dfm_1,
          sigmoid_table_965_0_sva_dfm_1, sigmoid_table_966_0_sva_dfm_1, sigmoid_table_967_0_sva_dfm_1,
          sigmoid_table_968_0_sva_dfm_1, sigmoid_table_969_0_sva_dfm_1, sigmoid_table_970_0_sva_dfm_1,
          sigmoid_table_971_0_sva_dfm_1, sigmoid_table_972_0_sva_dfm_1, sigmoid_table_973_0_sva_dfm_1,
          sigmoid_table_974_0_sva_dfm_1, sigmoid_table_975_0_sva_dfm_1, sigmoid_table_976_0_sva_dfm_1,
          sigmoid_table_977_0_sva_dfm_1, sigmoid_table_978_0_sva_dfm_1, sigmoid_table_979_0_sva_dfm_1,
          sigmoid_table_980_0_sva_dfm_1, sigmoid_table_981_0_sva_dfm_1, sigmoid_table_982_0_sva_dfm_1,
          sigmoid_table_983_0_sva_dfm_1, sigmoid_table_984_0_sva_dfm_1, sigmoid_table_985_0_sva_dfm_1,
          sigmoid_table_986_0_sva_dfm_1, sigmoid_table_987_0_sva_dfm_1, sigmoid_table_988_0_sva_dfm_1,
          sigmoid_table_989_0_sva_dfm_1, sigmoid_table_990_0_sva_dfm_1, sigmoid_table_991_0_sva_dfm_1,
          sigmoid_table_992_0_sva_dfm_1, sigmoid_table_993_0_sva_dfm_1, sigmoid_table_994_0_sva_dfm_1,
          sigmoid_table_995_0_sva_dfm_1, sigmoid_table_996_0_sva_dfm_1, sigmoid_table_997_0_sva_dfm_1,
          sigmoid_table_998_0_sva_dfm_1, sigmoid_table_999_0_sva_dfm_1, sigmoid_table_1000_0_sva_dfm_1,
          sigmoid_table_1001_0_sva_dfm_1, sigmoid_table_1002_0_sva_dfm_1, sigmoid_table_1003_0_sva_dfm_1,
          sigmoid_table_1004_0_sva_dfm_1, sigmoid_table_1005_0_sva_dfm_1, sigmoid_table_1006_0_sva_dfm_1,
          sigmoid_table_1007_0_sva_dfm_1, sigmoid_table_1008_0_sva_dfm_1, sigmoid_table_1009_0_sva_dfm_1,
          sigmoid_table_1010_0_sva_dfm_1, sigmoid_table_1011_0_sva_dfm_1, sigmoid_table_1012_0_sva_dfm_1,
          sigmoid_table_1013_0_sva_dfm_1, sigmoid_table_1014_0_sva_dfm_1, sigmoid_table_1015_0_sva_dfm_1,
          sigmoid_table_1016_0_sva_dfm_1, sigmoid_table_1017_0_sva_dfm_1, sigmoid_table_1018_0_sva_dfm_1,
          sigmoid_table_1019_0_sva_dfm_1, sigmoid_table_1020_0_sva_dfm_1, sigmoid_table_1021_0_sva_dfm_1,
          sigmoid_table_1022_0_sva_dfm_1, sigmoid_table_1023_0_sva_dfm_1, {for_for_or_1_itm
          , for_for_or_itm});
      res_rsci_d_1 <= MUX_s_1_1024_2(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_113_1_sva_dfm_1,
          sigmoid_table_114_1_sva_dfm_1, sigmoid_table_115_1_sva_dfm_1, sigmoid_table_116_1_sva_dfm_1,
          sigmoid_table_117_1_sva_dfm_1, sigmoid_table_118_1_sva_dfm_1, sigmoid_table_119_1_sva_dfm_1,
          sigmoid_table_120_1_sva_dfm_1, sigmoid_table_121_1_sva_dfm_1, sigmoid_table_122_1_sva_dfm_1,
          sigmoid_table_123_1_sva_dfm_1, sigmoid_table_124_1_sva_dfm_1, sigmoid_table_125_1_sva_dfm_1,
          sigmoid_table_126_1_sva_dfm_1, sigmoid_table_127_1_sva_dfm_1, sigmoid_table_128_1_sva_dfm_1,
          sigmoid_table_129_1_sva_dfm_1, sigmoid_table_130_1_sva_dfm_1, sigmoid_table_131_1_sva_dfm_1,
          sigmoid_table_132_1_sva_dfm_1, sigmoid_table_133_1_sva_dfm_1, sigmoid_table_134_1_sva_dfm_1,
          sigmoid_table_135_1_sva_dfm_1, sigmoid_table_136_1_sva_dfm_1, sigmoid_table_137_1_sva_dfm_1,
          sigmoid_table_138_1_sva_dfm_1, sigmoid_table_139_0_sva_dfm_1, sigmoid_table_140_0_sva_dfm_1,
          sigmoid_table_141_0_sva_dfm_1, sigmoid_table_142_0_sva_dfm_1, sigmoid_table_143_0_sva_dfm_1,
          sigmoid_table_144_0_sva_dfm_1, sigmoid_table_145_0_sva_dfm_1, sigmoid_table_146_0_sva_dfm_1,
          sigmoid_table_147_0_sva_dfm_1, sigmoid_table_148_0_sva_dfm_1, sigmoid_table_149_0_sva_dfm_1,
          sigmoid_table_150_0_sva_dfm_1, sigmoid_table_151_0_sva_dfm_1, sigmoid_table_152_0_sva_dfm_1,
          sigmoid_table_153_0_sva_dfm_1, sigmoid_table_154_0_sva_dfm_1, sigmoid_table_155_0_sva_dfm_1,
          sigmoid_table_156_0_sva_dfm_1, sigmoid_table_157_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          sigmoid_table_184_1_sva_dfm_1, sigmoid_table_185_1_sva_dfm_1, sigmoid_table_186_1_sva_dfm_1,
          sigmoid_table_187_1_sva_dfm_1, sigmoid_table_188_1_sva_dfm_1, sigmoid_table_189_1_sva_dfm_1,
          sigmoid_table_190_1_sva_dfm_1, sigmoid_table_191_1_sva_dfm_1, sigmoid_table_192_1_sva_dfm_1,
          sigmoid_table_193_1_sva_dfm_1, sigmoid_table_194_0_sva_dfm_1, sigmoid_table_195_0_sva_dfm_1,
          sigmoid_table_196_0_sva_dfm_1, sigmoid_table_197_0_sva_dfm_1, sigmoid_table_198_0_sva_dfm_1,
          sigmoid_table_199_0_sva_dfm_1, sigmoid_table_200_0_sva_dfm_1, sigmoid_table_201_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, sigmoid_table_217_1_sva_dfm_1, sigmoid_table_218_1_sva_dfm_1,
          sigmoid_table_219_1_sva_dfm_1, sigmoid_table_220_1_sva_dfm_1, sigmoid_table_221_1_sva_dfm_1,
          sigmoid_table_222_1_sva_dfm_1, sigmoid_table_223_0_sva_dfm_1, sigmoid_table_224_0_sva_dfm_1,
          sigmoid_table_225_0_sva_dfm_1, sigmoid_table_226_0_sva_dfm_1, sigmoid_table_227_0_sva_dfm_1,
          sigmoid_table_228_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, sigmoid_table_239_1_sva_dfm_1, sigmoid_table_240_1_sva_dfm_1,
          sigmoid_table_241_1_sva_dfm_1, sigmoid_table_242_1_sva_dfm_1, sigmoid_table_243_0_sva_dfm_1,
          sigmoid_table_244_0_sva_dfm_1, sigmoid_table_245_0_sva_dfm_1, sigmoid_table_246_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_255_1_sva_dfm_1,
          sigmoid_table_256_1_sva_dfm_1, sigmoid_table_257_1_sva_dfm_1, sigmoid_table_258_1_sva_dfm_1,
          sigmoid_table_259_0_sva_dfm_1, sigmoid_table_260_0_sva_dfm_1, sigmoid_table_261_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_268_1_sva_dfm_1, sigmoid_table_269_1_sva_dfm_1,
          sigmoid_table_270_1_sva_dfm_1, sigmoid_table_271_0_sva_dfm_1, sigmoid_table_272_0_sva_dfm_1,
          sigmoid_table_273_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_279_1_sva_dfm_1,
          sigmoid_table_280_1_sva_dfm_1, sigmoid_table_281_1_sva_dfm_1, sigmoid_table_282_0_sva_dfm_1,
          sigmoid_table_283_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_288_1_sva_dfm_1,
          sigmoid_table_289_1_sva_dfm_1, sigmoid_table_290_1_sva_dfm_1, sigmoid_table_291_0_sva_dfm_1,
          sigmoid_table_292_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_297_1_sva_dfm_1,
          sigmoid_table_298_1_sva_dfm_1, sigmoid_table_299_0_sva_dfm_1, sigmoid_table_300_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, sigmoid_table_304_1_sva_dfm_1, sigmoid_table_305_1_sva_dfm_1,
          sigmoid_table_306_0_sva_dfm_1, sigmoid_table_307_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, sigmoid_table_311_1_sva_dfm_1, sigmoid_table_312_0_sva_dfm_1, sigmoid_table_313_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, sigmoid_table_317_1_sva_dfm_1, sigmoid_table_318_0_sva_dfm_1,
          sigmoid_table_319_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_322_1_sva_dfm_1,
          sigmoid_table_323_1_sva_dfm_1, sigmoid_table_324_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, sigmoid_table_328_1_sva_dfm_1, sigmoid_table_329_0_sva_dfm_1, 1'b0,
          1'b0, sigmoid_table_332_1_sva_dfm_1, sigmoid_table_333_1_sva_dfm_1, sigmoid_table_334_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_337_1_sva_dfm_1, sigmoid_table_338_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_341_1_sva_dfm_1, sigmoid_table_342_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_345_1_sva_dfm_1, sigmoid_table_346_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_349_1_sva_dfm_1, sigmoid_table_350_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_353_1_sva_dfm_1, sigmoid_table_354_0_sva_dfm_1,
          1'b0, sigmoid_table_356_1_sva_dfm_1, sigmoid_table_357_0_sva_dfm_1, 1'b0,
          1'b0, sigmoid_table_360_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_363_1_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_366_1_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_369_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_372_0_sva_dfm_1, 1'b0, sigmoid_table_374_1_sva_dfm_1,
          sigmoid_table_375_0_sva_dfm_1, 1'b0, sigmoid_table_377_1_sva_dfm_1, 1'b0,
          1'b0, sigmoid_table_380_0_sva_dfm_1, 1'b0, sigmoid_table_382_1_sva_dfm_1,
          1'b0, sigmoid_table_384_1_sva_dfm_1, sigmoid_table_385_0_sva_dfm_1, 1'b0,
          sigmoid_table_387_0_sva_dfm_1, 1'b0, sigmoid_table_389_1_sva_dfm_1, 1'b0,
          sigmoid_table_391_1_sva_dfm_1, 1'b0, sigmoid_table_393_1_sva_dfm_1, sigmoid_table_394_0_sva_dfm_1,
          1'b0, sigmoid_table_396_0_sva_dfm_1, 1'b0, sigmoid_table_398_0_sva_dfm_1,
          1'b0, sigmoid_table_400_0_sva_dfm_1, 1'b0, sigmoid_table_402_0_sva_dfm_1,
          1'b0, sigmoid_table_404_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_407_1_sva_dfm_1,
          1'b0, sigmoid_table_409_1_sva_dfm_1, 1'b0, sigmoid_table_411_0_sva_dfm_1,
          1'b0, sigmoid_table_413_0_sva_dfm_1, sigmoid_table_414_1_sva_dfm_1, 1'b0,
          sigmoid_table_416_1_sva_dfm_1, 1'b0, sigmoid_table_418_0_sva_dfm_1, sigmoid_table_419_1_sva_dfm_1,
          1'b0, sigmoid_table_421_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_424_1_sva_dfm_1,
          1'b0, sigmoid_table_426_0_sva_dfm_1, sigmoid_table_427_1_sva_dfm_1, 1'b0,
          sigmoid_table_429_0_sva_dfm_1, sigmoid_table_430_1_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_433_1_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_436_0_sva_dfm_1,
          sigmoid_table_437_1_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_440_1_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_443_0_sva_dfm_1, sigmoid_table_444_1_sva_dfm_1,
          sigmoid_table_445_1_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_448_0_sva_dfm_1,
          sigmoid_table_449_1_sva_dfm_1, 1'b0, 1'b0, 1'b0, sigmoid_table_453_0_sva_dfm_1,
          sigmoid_table_454_1_sva_dfm_1, 1'b0, 1'b0, 1'b0, sigmoid_table_458_0_sva_dfm_1,
          sigmoid_table_459_0_sva_dfm_1, sigmoid_table_460_1_sva_dfm_1, sigmoid_table_461_1_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_466_0_sva_dfm_1, sigmoid_table_467_0_sva_dfm_1,
          sigmoid_table_468_1_sva_dfm_1, sigmoid_table_469_1_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, sigmoid_table_475_0_sva_dfm_1, sigmoid_table_476_0_sva_dfm_1,
          sigmoid_table_477_0_sva_dfm_1, sigmoid_table_478_0_sva_dfm_1, sigmoid_table_479_1_sva_dfm_1,
          sigmoid_table_480_1_sva_dfm_1, sigmoid_table_481_1_sva_dfm_1, sigmoid_table_482_1_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_516_0_sva_dfm_1,
          sigmoid_table_517_0_sva_dfm_1, sigmoid_table_518_0_sva_dfm_1, sigmoid_table_519_0_sva_dfm_1,
          sigmoid_table_520_0_sva_dfm_1, sigmoid_table_521_0_sva_dfm_1, sigmoid_table_522_0_sva_dfm_1,
          sigmoid_table_523_0_sva_dfm_1, sigmoid_table_524_0_sva_dfm_1, sigmoid_table_525_0_sva_dfm_1,
          sigmoid_table_526_0_sva_dfm_1, sigmoid_table_527_0_sva_dfm_1, sigmoid_table_528_0_sva_dfm_1,
          sigmoid_table_529_0_sva_dfm_1, sigmoid_table_530_0_sva_dfm_1, sigmoid_table_531_0_sva_dfm_1,
          sigmoid_table_532_0_sva_dfm_1, sigmoid_table_533_0_sva_dfm_1, sigmoid_table_534_0_sva_dfm_1,
          sigmoid_table_535_0_sva_dfm_1, sigmoid_table_536_1_sva_dfm_1, sigmoid_table_537_1_sva_dfm_1,
          sigmoid_table_538_1_sva_dfm_1, sigmoid_table_539_1_sva_dfm_1, sigmoid_table_540_1_sva_dfm_1,
          sigmoid_table_541_1_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, sigmoid_table_550_0_sva_dfm_1, sigmoid_table_551_0_sva_dfm_1, sigmoid_table_552_1_sva_dfm_1,
          sigmoid_table_553_1_sva_dfm_1, sigmoid_table_554_1_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_559_0_sva_dfm_1, sigmoid_table_560_0_sva_dfm_1,
          sigmoid_table_561_1_sva_dfm_1, sigmoid_table_562_1_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_567_0_sva_dfm_1, sigmoid_table_568_1_sva_dfm_1,
          sigmoid_table_569_1_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_572_0_sva_dfm_1,
          sigmoid_table_573_0_sva_dfm_1, sigmoid_table_574_1_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_577_0_sva_dfm_1, sigmoid_table_578_1_sva_dfm_1, 1'b0, 1'b0,
          1'b0, sigmoid_table_582_0_sva_dfm_1, sigmoid_table_583_1_sva_dfm_1, 1'b0,
          sigmoid_table_585_0_sva_dfm_1, sigmoid_table_586_1_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_589_0_sva_dfm_1, sigmoid_table_590_1_sva_dfm_1, 1'b0, sigmoid_table_592_0_sva_dfm_1,
          sigmoid_table_593_1_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_596_1_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_599_1_sva_dfm_1, 1'b0, sigmoid_table_601_0_sva_dfm_1,
          sigmoid_table_602_1_sva_dfm_1, 1'b0, sigmoid_table_604_0_sva_dfm_1, 1'b0,
          1'b0, sigmoid_table_607_1_sva_dfm_1, 1'b0, sigmoid_table_609_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_612_1_sva_dfm_1, 1'b0, sigmoid_table_614_0_sva_dfm_1,
          1'b0, sigmoid_table_616_0_sva_dfm_1, 1'b0, sigmoid_table_618_0_sva_dfm_1,
          sigmoid_table_619_1_sva_dfm_1, 1'b0, sigmoid_table_621_1_sva_dfm_1, 1'b0,
          sigmoid_table_623_1_sva_dfm_1, 1'b0, sigmoid_table_625_1_sva_dfm_1, 1'b0,
          sigmoid_table_627_1_sva_dfm_1, 1'b0, sigmoid_table_629_1_sva_dfm_1, 1'b0,
          1'b0, sigmoid_table_632_0_sva_dfm_1, 1'b0, sigmoid_table_634_0_sva_dfm_1,
          1'b0, sigmoid_table_636_0_sva_dfm_1, 1'b0, sigmoid_table_638_1_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_641_0_sva_dfm_1, 1'b0, sigmoid_table_643_1_sva_dfm_1,
          1'b0, sigmoid_table_645_1_sva_dfm_1, sigmoid_table_646_0_sva_dfm_1, 1'b0,
          sigmoid_table_648_1_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_651_0_sva_dfm_1,
          1'b0, sigmoid_table_653_1_sva_dfm_1, sigmoid_table_654_0_sva_dfm_1, 1'b0,
          sigmoid_table_656_1_sva_dfm_1, sigmoid_table_657_0_sva_dfm_1, 1'b0, sigmoid_table_659_1_sva_dfm_1,
          sigmoid_table_660_0_sva_dfm_1, 1'b0, sigmoid_table_662_1_sva_dfm_1, sigmoid_table_663_0_sva_dfm_1,
          1'b0, sigmoid_table_665_1_sva_dfm_1, sigmoid_table_666_0_sva_dfm_1, 1'b0,
          1'b0, sigmoid_table_669_1_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_672_1_sva_dfm_1,
          sigmoid_table_673_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_676_1_sva_dfm_1,
          sigmoid_table_677_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_680_1_sva_dfm_1,
          sigmoid_table_681_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_684_1_sva_dfm_1,
          sigmoid_table_685_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_688_1_sva_dfm_1,
          sigmoid_table_689_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, sigmoid_table_693_1_sva_dfm_1,
          sigmoid_table_694_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_697_1_sva_dfm_1,
          sigmoid_table_698_1_sva_dfm_1, sigmoid_table_699_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, sigmoid_table_703_1_sva_dfm_1, sigmoid_table_704_0_sva_dfm_1, 1'b0,
          1'b0, 1'b0, sigmoid_table_708_1_sva_dfm_1, sigmoid_table_709_1_sva_dfm_1,
          sigmoid_table_710_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, sigmoid_table_714_1_sva_dfm_1,
          sigmoid_table_715_1_sva_dfm_1, sigmoid_table_716_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_721_1_sva_dfm_1, sigmoid_table_722_1_sva_dfm_1,
          sigmoid_table_723_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_728_1_sva_dfm_1,
          sigmoid_table_729_1_sva_dfm_1, sigmoid_table_730_0_sva_dfm_1, sigmoid_table_731_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_737_1_sva_dfm_1, sigmoid_table_738_1_sva_dfm_1,
          sigmoid_table_739_0_sva_dfm_1, sigmoid_table_740_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, sigmoid_table_746_1_sva_dfm_1, sigmoid_table_747_1_sva_dfm_1,
          sigmoid_table_748_0_sva_dfm_1, sigmoid_table_749_0_sva_dfm_1, sigmoid_table_750_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_757_1_sva_dfm_1, sigmoid_table_758_1_sva_dfm_1,
          sigmoid_table_759_1_sva_dfm_1, sigmoid_table_760_0_sva_dfm_1, sigmoid_table_761_0_sva_dfm_1,
          sigmoid_table_762_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          sigmoid_table_770_1_sva_dfm_1, sigmoid_table_771_1_sva_dfm_1, sigmoid_table_772_1_sva_dfm_1,
          sigmoid_table_773_1_sva_dfm_1, sigmoid_table_774_0_sva_dfm_1, sigmoid_table_775_0_sva_dfm_1,
          sigmoid_table_776_0_sva_dfm_1, sigmoid_table_777_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_786_1_sva_dfm_1, sigmoid_table_787_1_sva_dfm_1,
          sigmoid_table_788_1_sva_dfm_1, sigmoid_table_789_1_sva_dfm_1, sigmoid_table_790_1_sva_dfm_1,
          sigmoid_table_791_0_sva_dfm_1, sigmoid_table_792_0_sva_dfm_1, sigmoid_table_793_0_sva_dfm_1,
          sigmoid_table_794_0_sva_dfm_1, sigmoid_table_795_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_808_1_sva_dfm_1,
          sigmoid_table_809_1_sva_dfm_1, sigmoid_table_810_1_sva_dfm_1, sigmoid_table_811_1_sva_dfm_1,
          sigmoid_table_812_1_sva_dfm_1, sigmoid_table_813_1_sva_dfm_1, sigmoid_table_814_1_sva_dfm_1,
          sigmoid_table_815_0_sva_dfm_1, sigmoid_table_816_0_sva_dfm_1, sigmoid_table_817_0_sva_dfm_1,
          sigmoid_table_818_0_sva_dfm_1, sigmoid_table_819_0_sva_dfm_1, sigmoid_table_820_0_sva_dfm_1,
          sigmoid_table_821_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          sigmoid_table_841_1_sva_dfm_1, sigmoid_table_842_1_sva_dfm_1, sigmoid_table_843_1_sva_dfm_1,
          sigmoid_table_844_1_sva_dfm_1, sigmoid_table_845_1_sva_dfm_1, sigmoid_table_846_1_sva_dfm_1,
          sigmoid_table_847_1_sva_dfm_1, sigmoid_table_848_1_sva_dfm_1, sigmoid_table_849_1_sva_dfm_1,
          sigmoid_table_850_1_sva_dfm_1, sigmoid_table_851_1_sva_dfm_1, sigmoid_table_852_1_sva_dfm_1,
          sigmoid_table_853_0_sva_dfm_1, sigmoid_table_854_0_sva_dfm_1, sigmoid_table_855_0_sva_dfm_1,
          sigmoid_table_856_0_sva_dfm_1, sigmoid_table_857_0_sva_dfm_1, sigmoid_table_858_0_sva_dfm_1,
          sigmoid_table_859_0_sva_dfm_1, sigmoid_table_860_0_sva_dfm_1, sigmoid_table_861_0_sva_dfm_1,
          sigmoid_table_862_0_sva_dfm_1, sigmoid_table_863_0_sva_dfm_1, sigmoid_table_864_0_sva_dfm_1,
          sigmoid_table_865_0_sva_dfm_1, sigmoid_table_866_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_911_1_sva_dfm_1, sigmoid_table_912_1_sva_dfm_1,
          sigmoid_table_913_1_sva_dfm_1, sigmoid_table_914_1_sva_dfm_1, sigmoid_table_915_1_sva_dfm_1,
          sigmoid_table_916_1_sva_dfm_1, sigmoid_table_917_1_sva_dfm_1, sigmoid_table_918_1_sva_dfm_1,
          sigmoid_table_919_1_sva_dfm_1, sigmoid_table_920_1_sva_dfm_1, sigmoid_table_921_1_sva_dfm_1,
          sigmoid_table_922_1_sva_dfm_1, sigmoid_table_923_1_sva_dfm_1, sigmoid_table_924_1_sva_dfm_1,
          sigmoid_table_925_1_sva_dfm_1, sigmoid_table_926_1_sva_dfm_1, sigmoid_table_927_1_sva_dfm_1,
          sigmoid_table_928_1_sva_dfm_1, sigmoid_table_929_1_sva_dfm_1, sigmoid_table_930_1_sva_dfm_1,
          sigmoid_table_931_1_sva_dfm_1, sigmoid_table_932_1_sva_dfm_1, sigmoid_table_933_1_sva_dfm_1,
          sigmoid_table_934_1_sva_dfm_1, sigmoid_table_935_1_sva_dfm_1, sigmoid_table_936_1_sva_dfm_1,
          sigmoid_table_937_1_sva_dfm_1, sigmoid_table_938_1_sva_dfm_1, sigmoid_table_939_1_sva_dfm_1,
          sigmoid_table_940_1_sva_dfm_1, sigmoid_table_941_1_sva_dfm_1, sigmoid_table_942_1_sva_dfm_1,
          sigmoid_table_943_1_sva_dfm_1, sigmoid_table_944_1_sva_dfm_1, sigmoid_table_945_1_sva_dfm_1,
          sigmoid_table_946_1_sva_dfm_1, sigmoid_table_947_1_sva_dfm_1, sigmoid_table_948_1_sva_dfm_1,
          sigmoid_table_949_1_sva_dfm_1, sigmoid_table_950_1_sva_dfm_1, sigmoid_table_951_1_sva_dfm_1,
          sigmoid_table_952_1_sva_dfm_1, sigmoid_table_953_1_sva_dfm_1, sigmoid_table_954_1_sva_dfm_1,
          sigmoid_table_955_0_sva_dfm_1, sigmoid_table_956_0_sva_dfm_1, sigmoid_table_957_0_sva_dfm_1,
          sigmoid_table_958_0_sva_dfm_1, sigmoid_table_959_0_sva_dfm_1, sigmoid_table_960_0_sva_dfm_1,
          sigmoid_table_961_0_sva_dfm_1, sigmoid_table_962_0_sva_dfm_1, sigmoid_table_963_0_sva_dfm_1,
          sigmoid_table_964_0_sva_dfm_1, sigmoid_table_965_0_sva_dfm_1, sigmoid_table_966_0_sva_dfm_1,
          sigmoid_table_967_0_sva_dfm_1, sigmoid_table_968_0_sva_dfm_1, sigmoid_table_969_0_sva_dfm_1,
          sigmoid_table_970_0_sva_dfm_1, sigmoid_table_971_0_sva_dfm_1, sigmoid_table_972_0_sva_dfm_1,
          sigmoid_table_973_0_sva_dfm_1, sigmoid_table_974_0_sva_dfm_1, sigmoid_table_975_0_sva_dfm_1,
          sigmoid_table_976_0_sva_dfm_1, sigmoid_table_977_0_sva_dfm_1, sigmoid_table_978_0_sva_dfm_1,
          sigmoid_table_979_0_sva_dfm_1, sigmoid_table_980_0_sva_dfm_1, sigmoid_table_981_0_sva_dfm_1,
          sigmoid_table_982_0_sva_dfm_1, sigmoid_table_983_0_sva_dfm_1, sigmoid_table_984_0_sva_dfm_1,
          sigmoid_table_985_0_sva_dfm_1, sigmoid_table_986_0_sva_dfm_1, sigmoid_table_987_0_sva_dfm_1,
          sigmoid_table_988_0_sva_dfm_1, sigmoid_table_989_0_sva_dfm_1, sigmoid_table_990_0_sva_dfm_1,
          sigmoid_table_991_0_sva_dfm_1, sigmoid_table_992_0_sva_dfm_1, sigmoid_table_993_0_sva_dfm_1,
          sigmoid_table_994_0_sva_dfm_1, sigmoid_table_995_0_sva_dfm_1, sigmoid_table_996_0_sva_dfm_1,
          sigmoid_table_997_0_sva_dfm_1, sigmoid_table_998_0_sva_dfm_1, sigmoid_table_999_0_sva_dfm_1,
          sigmoid_table_1000_0_sva_dfm_1, sigmoid_table_1001_0_sva_dfm_1, sigmoid_table_1002_0_sva_dfm_1,
          sigmoid_table_1003_0_sva_dfm_1, sigmoid_table_1004_0_sva_dfm_1, sigmoid_table_1005_0_sva_dfm_1,
          sigmoid_table_1006_0_sva_dfm_1, sigmoid_table_1007_0_sva_dfm_1, sigmoid_table_1008_0_sva_dfm_1,
          sigmoid_table_1009_0_sva_dfm_1, sigmoid_table_1010_0_sva_dfm_1, sigmoid_table_1011_0_sva_dfm_1,
          sigmoid_table_1012_0_sva_dfm_1, sigmoid_table_1013_0_sva_dfm_1, sigmoid_table_1014_0_sva_dfm_1,
          sigmoid_table_1015_0_sva_dfm_1, sigmoid_table_1016_0_sva_dfm_1, sigmoid_table_1017_0_sva_dfm_1,
          sigmoid_table_1018_0_sva_dfm_1, sigmoid_table_1019_0_sva_dfm_1, sigmoid_table_1020_0_sva_dfm_1,
          sigmoid_table_1021_0_sva_dfm_1, sigmoid_table_1022_0_sva_dfm_1, sigmoid_table_1023_0_sva_dfm_1,
          {for_for_or_1_itm , for_for_or_itm});
      res_rsci_d_8 <= MUX_s_1_1024_2(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_442_8_sva_dfm_1, sigmoid_table_443_8_sva_dfm_1,
          sigmoid_table_444_8_sva_dfm_1, sigmoid_table_445_8_sva_dfm_1, sigmoid_table_446_8_sva_dfm_1,
          sigmoid_table_447_8_sva_dfm_1, sigmoid_table_448_8_sva_dfm_1, sigmoid_table_449_8_sva_dfm_1,
          sigmoid_table_450_8_sva_dfm_1, sigmoid_table_451_8_sva_dfm_1, sigmoid_table_452_8_sva_dfm_1,
          sigmoid_table_453_8_sva_dfm_1, sigmoid_table_454_8_sva_dfm_1, sigmoid_table_455_8_sva_dfm_1,
          sigmoid_table_456_8_sva_dfm_1, sigmoid_table_457_8_sva_dfm_1, sigmoid_table_458_8_sva_dfm_1,
          sigmoid_table_459_8_sva_dfm_1, sigmoid_table_460_8_sva_dfm_1, sigmoid_table_461_8_sva_dfm_1,
          sigmoid_table_462_8_sva_dfm_1, sigmoid_table_463_8_sva_dfm_1, sigmoid_table_464_8_sva_dfm_1,
          sigmoid_table_465_8_sva_dfm_1, sigmoid_table_466_8_sva_dfm_1, sigmoid_table_467_8_sva_dfm_1,
          sigmoid_table_468_8_sva_dfm_1, sigmoid_table_469_8_sva_dfm_1, sigmoid_table_470_8_sva_dfm_1,
          sigmoid_table_471_8_sva_dfm_1, sigmoid_table_472_8_sva_dfm_1, sigmoid_table_473_8_sva_dfm_1,
          sigmoid_table_474_8_sva_dfm_1, sigmoid_table_475_8_sva_dfm_1, sigmoid_table_476_8_sva_dfm_1,
          sigmoid_table_477_8_sva_dfm_1, sigmoid_table_478_8_sva_dfm_1, sigmoid_table_479_8_sva_dfm_1,
          sigmoid_table_480_7_sva_dfm_1, sigmoid_table_481_7_sva_dfm_1, sigmoid_table_482_7_sva_dfm_1,
          sigmoid_table_483_7_sva_dfm_1, sigmoid_table_484_7_sva_dfm_1, sigmoid_table_485_7_sva_dfm_1,
          sigmoid_table_486_7_sva_dfm_1, sigmoid_table_487_7_sva_dfm_1, sigmoid_table_488_7_sva_dfm_1,
          sigmoid_table_489_7_sva_dfm_1, sigmoid_table_490_7_sva_dfm_1, sigmoid_table_491_7_sva_dfm_1,
          sigmoid_table_492_7_sva_dfm_1, sigmoid_table_493_7_sva_dfm_1, sigmoid_table_494_7_sva_dfm_1,
          sigmoid_table_495_7_sva_dfm_1, sigmoid_table_496_6_sva_dfm_1, sigmoid_table_497_6_sva_dfm_1,
          sigmoid_table_498_6_sva_dfm_1, sigmoid_table_499_6_sva_dfm_1, sigmoid_table_500_6_sva_dfm_1,
          sigmoid_table_501_6_sva_dfm_1, sigmoid_table_502_6_sva_dfm_1, sigmoid_table_503_6_sva_dfm_1,
          sigmoid_table_504_5_sva_dfm_1, sigmoid_table_505_5_sva_dfm_1, sigmoid_table_506_5_sva_dfm_1,
          sigmoid_table_507_5_sva_dfm_1, sigmoid_table_508_4_sva_dfm_1, sigmoid_table_509_4_sva_dfm_1,
          sigmoid_table_510_3_sva_dfm_1, sigmoid_table_511_2_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_583_8_sva_dfm_1,
          sigmoid_table_584_8_sva_dfm_1, sigmoid_table_585_8_sva_dfm_1, sigmoid_table_586_8_sva_dfm_1,
          sigmoid_table_587_8_sva_dfm_1, sigmoid_table_588_8_sva_dfm_1, sigmoid_table_589_8_sva_dfm_1,
          sigmoid_table_590_8_sva_dfm_1, sigmoid_table_591_8_sva_dfm_1, sigmoid_table_592_8_sva_dfm_1,
          sigmoid_table_593_8_sva_dfm_1, sigmoid_table_594_8_sva_dfm_1, sigmoid_table_595_8_sva_dfm_1,
          sigmoid_table_596_8_sva_dfm_1, sigmoid_table_597_8_sva_dfm_1, sigmoid_table_598_8_sva_dfm_1,
          sigmoid_table_599_8_sva_dfm_1, sigmoid_table_600_8_sva_dfm_1, sigmoid_table_601_8_sva_dfm_1,
          sigmoid_table_602_8_sva_dfm_1, sigmoid_table_603_8_sva_dfm_1, sigmoid_table_604_8_sva_dfm_1,
          sigmoid_table_605_8_sva_dfm_1, sigmoid_table_606_8_sva_dfm_1, sigmoid_table_607_8_sva_dfm_1,
          sigmoid_table_608_8_sva_dfm_1, sigmoid_table_609_8_sva_dfm_1, sigmoid_table_610_8_sva_dfm_1,
          sigmoid_table_611_8_sva_dfm_1, sigmoid_table_612_8_sva_dfm_1, sigmoid_table_613_8_sva_dfm_1,
          sigmoid_table_614_8_sva_dfm_1, sigmoid_table_615_8_sva_dfm_1, sigmoid_table_616_8_sva_dfm_1,
          sigmoid_table_617_8_sva_dfm_1, sigmoid_table_618_8_sva_dfm_1, sigmoid_table_619_8_sva_dfm_1,
          sigmoid_table_620_8_sva_dfm_1, sigmoid_table_621_8_sva_dfm_1, sigmoid_table_622_8_sva_dfm_1,
          sigmoid_table_623_8_sva_dfm_1, sigmoid_table_624_8_sva_dfm_1, sigmoid_table_625_8_sva_dfm_1,
          sigmoid_table_626_8_sva_dfm_1, sigmoid_table_627_8_sva_dfm_1, sigmoid_table_628_8_sva_dfm_1,
          sigmoid_table_629_8_sva_dfm_1, sigmoid_table_630_8_sva_dfm_1, sigmoid_table_631_8_sva_dfm_1,
          sigmoid_table_632_8_sva_dfm_1, sigmoid_table_633_8_sva_dfm_1, sigmoid_table_634_8_sva_dfm_1,
          sigmoid_table_635_8_sva_dfm_1, sigmoid_table_636_8_sva_dfm_1, sigmoid_table_637_7_sva_dfm_1,
          sigmoid_table_638_7_sva_dfm_1, sigmoid_table_639_7_sva_dfm_1, sigmoid_table_640_7_sva_dfm_1,
          sigmoid_table_641_7_sva_dfm_1, sigmoid_table_642_7_sva_dfm_1, sigmoid_table_643_7_sva_dfm_1,
          sigmoid_table_644_7_sva_dfm_1, sigmoid_table_645_7_sva_dfm_1, sigmoid_table_646_7_sva_dfm_1,
          sigmoid_table_647_7_sva_dfm_1, sigmoid_table_648_7_sva_dfm_1, sigmoid_table_649_7_sva_dfm_1,
          sigmoid_table_650_7_sva_dfm_1, sigmoid_table_651_7_sva_dfm_1, sigmoid_table_652_7_sva_dfm_1,
          sigmoid_table_653_7_sva_dfm_1, sigmoid_table_654_7_sva_dfm_1, sigmoid_table_655_7_sva_dfm_1,
          sigmoid_table_656_7_sva_dfm_1, sigmoid_table_657_7_sva_dfm_1, sigmoid_table_658_7_sva_dfm_1,
          sigmoid_table_659_7_sva_dfm_1, sigmoid_table_660_7_sva_dfm_1, sigmoid_table_661_7_sva_dfm_1,
          sigmoid_table_662_7_sva_dfm_1, sigmoid_table_663_7_sva_dfm_1, sigmoid_table_664_7_sva_dfm_1,
          sigmoid_table_665_7_sva_dfm_1, sigmoid_table_666_7_sva_dfm_1, sigmoid_table_667_7_sva_dfm_1,
          sigmoid_table_668_7_sva_dfm_1, sigmoid_table_669_7_sva_dfm_1, sigmoid_table_670_7_sva_dfm_1,
          sigmoid_table_671_7_sva_dfm_1, sigmoid_table_672_7_sva_dfm_1, sigmoid_table_673_7_sva_dfm_1,
          sigmoid_table_674_7_sva_dfm_1, sigmoid_table_675_7_sva_dfm_1, sigmoid_table_676_7_sva_dfm_1,
          sigmoid_table_677_7_sva_dfm_1, sigmoid_table_678_7_sva_dfm_1, sigmoid_table_679_7_sva_dfm_1,
          sigmoid_table_680_7_sva_dfm_1, sigmoid_table_681_7_sva_dfm_1, sigmoid_table_682_7_sva_dfm_1,
          sigmoid_table_683_7_sva_dfm_1, sigmoid_table_684_7_sva_dfm_1, sigmoid_table_685_7_sva_dfm_1,
          sigmoid_table_686_6_sva_dfm_1, sigmoid_table_687_6_sva_dfm_1, sigmoid_table_688_6_sva_dfm_1,
          sigmoid_table_689_6_sva_dfm_1, sigmoid_table_690_6_sva_dfm_1, sigmoid_table_691_6_sva_dfm_1,
          sigmoid_table_692_6_sva_dfm_1, sigmoid_table_693_6_sva_dfm_1, sigmoid_table_694_6_sva_dfm_1,
          sigmoid_table_695_6_sva_dfm_1, sigmoid_table_696_6_sva_dfm_1, sigmoid_table_697_6_sva_dfm_1,
          sigmoid_table_698_6_sva_dfm_1, sigmoid_table_699_6_sva_dfm_1, sigmoid_table_700_6_sva_dfm_1,
          sigmoid_table_701_6_sva_dfm_1, sigmoid_table_702_6_sva_dfm_1, sigmoid_table_703_6_sva_dfm_1,
          sigmoid_table_704_6_sva_dfm_1, sigmoid_table_705_6_sva_dfm_1, sigmoid_table_706_6_sva_dfm_1,
          sigmoid_table_707_6_sva_dfm_1, sigmoid_table_708_6_sva_dfm_1, sigmoid_table_709_6_sva_dfm_1,
          sigmoid_table_710_6_sva_dfm_1, sigmoid_table_711_6_sva_dfm_1, sigmoid_table_712_6_sva_dfm_1,
          sigmoid_table_713_6_sva_dfm_1, sigmoid_table_714_6_sva_dfm_1, sigmoid_table_715_6_sva_dfm_1,
          sigmoid_table_716_6_sva_dfm_1, sigmoid_table_717_6_sva_dfm_1, sigmoid_table_718_6_sva_dfm_1,
          sigmoid_table_719_6_sva_dfm_1, sigmoid_table_720_6_sva_dfm_1, sigmoid_table_721_6_sva_dfm_1,
          sigmoid_table_722_6_sva_dfm_1, sigmoid_table_723_6_sva_dfm_1, sigmoid_table_724_6_sva_dfm_1,
          sigmoid_table_725_6_sva_dfm_1, sigmoid_table_726_6_sva_dfm_1, sigmoid_table_727_6_sva_dfm_1,
          sigmoid_table_728_6_sva_dfm_1, sigmoid_table_729_6_sva_dfm_1, sigmoid_table_730_6_sva_dfm_1,
          sigmoid_table_731_6_sva_dfm_1, sigmoid_table_732_5_sva_dfm_1, sigmoid_table_733_5_sva_dfm_1,
          sigmoid_table_734_5_sva_dfm_1, sigmoid_table_735_5_sva_dfm_1, sigmoid_table_736_5_sva_dfm_1,
          sigmoid_table_737_5_sva_dfm_1, sigmoid_table_738_5_sva_dfm_1, sigmoid_table_739_5_sva_dfm_1,
          sigmoid_table_740_5_sva_dfm_1, sigmoid_table_741_5_sva_dfm_1, sigmoid_table_742_5_sva_dfm_1,
          sigmoid_table_743_5_sva_dfm_1, sigmoid_table_744_5_sva_dfm_1, sigmoid_table_745_5_sva_dfm_1,
          sigmoid_table_746_5_sva_dfm_1, sigmoid_table_747_5_sva_dfm_1, sigmoid_table_748_5_sva_dfm_1,
          sigmoid_table_749_5_sva_dfm_1, sigmoid_table_750_5_sva_dfm_1, sigmoid_table_751_5_sva_dfm_1,
          sigmoid_table_752_5_sva_dfm_1, sigmoid_table_753_5_sva_dfm_1, sigmoid_table_754_5_sva_dfm_1,
          sigmoid_table_755_5_sva_dfm_1, sigmoid_table_756_5_sva_dfm_1, sigmoid_table_757_5_sva_dfm_1,
          sigmoid_table_758_5_sva_dfm_1, sigmoid_table_759_5_sva_dfm_1, sigmoid_table_760_5_sva_dfm_1,
          sigmoid_table_761_5_sva_dfm_1, sigmoid_table_762_5_sva_dfm_1, sigmoid_table_763_5_sva_dfm_1,
          sigmoid_table_764_5_sva_dfm_1, sigmoid_table_765_5_sva_dfm_1, sigmoid_table_766_5_sva_dfm_1,
          sigmoid_table_767_5_sva_dfm_1, sigmoid_table_768_5_sva_dfm_1, sigmoid_table_769_5_sva_dfm_1,
          sigmoid_table_770_5_sva_dfm_1, sigmoid_table_771_5_sva_dfm_1, sigmoid_table_772_5_sva_dfm_1,
          sigmoid_table_773_5_sva_dfm_1, sigmoid_table_774_5_sva_dfm_1, sigmoid_table_775_5_sva_dfm_1,
          sigmoid_table_776_5_sva_dfm_1, sigmoid_table_777_5_sva_dfm_1, sigmoid_table_778_4_sva_dfm_1,
          sigmoid_table_779_4_sva_dfm_1, sigmoid_table_780_4_sva_dfm_1, sigmoid_table_781_4_sva_dfm_1,
          sigmoid_table_782_4_sva_dfm_1, sigmoid_table_783_4_sva_dfm_1, sigmoid_table_784_4_sva_dfm_1,
          sigmoid_table_785_4_sva_dfm_1, sigmoid_table_786_4_sva_dfm_1, sigmoid_table_787_4_sva_dfm_1,
          sigmoid_table_788_4_sva_dfm_1, sigmoid_table_789_4_sva_dfm_1, sigmoid_table_790_4_sva_dfm_1,
          sigmoid_table_791_4_sva_dfm_1, sigmoid_table_792_4_sva_dfm_1, sigmoid_table_793_4_sva_dfm_1,
          sigmoid_table_794_4_sva_dfm_1, sigmoid_table_795_4_sva_dfm_1, sigmoid_table_796_4_sva_dfm_1,
          sigmoid_table_797_4_sva_dfm_1, sigmoid_table_798_4_sva_dfm_1, sigmoid_table_799_4_sva_dfm_1,
          sigmoid_table_800_4_sva_dfm_1, sigmoid_table_801_4_sva_dfm_1, sigmoid_table_802_4_sva_dfm_1,
          sigmoid_table_803_4_sva_dfm_1, sigmoid_table_804_4_sva_dfm_1, sigmoid_table_805_4_sva_dfm_1,
          sigmoid_table_806_4_sva_dfm_1, sigmoid_table_807_4_sva_dfm_1, sigmoid_table_808_4_sva_dfm_1,
          sigmoid_table_809_4_sva_dfm_1, sigmoid_table_810_4_sva_dfm_1, sigmoid_table_811_4_sva_dfm_1,
          sigmoid_table_812_4_sva_dfm_1, sigmoid_table_813_4_sva_dfm_1, sigmoid_table_814_4_sva_dfm_1,
          sigmoid_table_815_4_sva_dfm_1, sigmoid_table_816_4_sva_dfm_1, sigmoid_table_817_4_sva_dfm_1,
          sigmoid_table_818_4_sva_dfm_1, sigmoid_table_819_4_sva_dfm_1, sigmoid_table_820_4_sva_dfm_1,
          sigmoid_table_821_4_sva_dfm_1, sigmoid_table_822_3_sva_dfm_1, sigmoid_table_823_3_sva_dfm_1,
          sigmoid_table_824_3_sva_dfm_1, sigmoid_table_825_3_sva_dfm_1, sigmoid_table_826_3_sva_dfm_1,
          sigmoid_table_827_3_sva_dfm_1, sigmoid_table_828_3_sva_dfm_1, sigmoid_table_829_3_sva_dfm_1,
          sigmoid_table_830_3_sva_dfm_1, sigmoid_table_831_3_sva_dfm_1, sigmoid_table_832_3_sva_dfm_1,
          sigmoid_table_833_3_sva_dfm_1, sigmoid_table_834_3_sva_dfm_1, sigmoid_table_835_3_sva_dfm_1,
          sigmoid_table_836_3_sva_dfm_1, sigmoid_table_837_3_sva_dfm_1, sigmoid_table_838_3_sva_dfm_1,
          sigmoid_table_839_3_sva_dfm_1, sigmoid_table_840_3_sva_dfm_1, sigmoid_table_841_3_sva_dfm_1,
          sigmoid_table_842_3_sva_dfm_1, sigmoid_table_843_3_sva_dfm_1, sigmoid_table_844_3_sva_dfm_1,
          sigmoid_table_845_3_sva_dfm_1, sigmoid_table_846_3_sva_dfm_1, sigmoid_table_847_3_sva_dfm_1,
          sigmoid_table_848_3_sva_dfm_1, sigmoid_table_849_3_sva_dfm_1, sigmoid_table_850_3_sva_dfm_1,
          sigmoid_table_851_3_sva_dfm_1, sigmoid_table_852_3_sva_dfm_1, sigmoid_table_853_3_sva_dfm_1,
          sigmoid_table_854_3_sva_dfm_1, sigmoid_table_855_3_sva_dfm_1, sigmoid_table_856_3_sva_dfm_1,
          sigmoid_table_857_3_sva_dfm_1, sigmoid_table_858_3_sva_dfm_1, sigmoid_table_859_3_sva_dfm_1,
          sigmoid_table_860_3_sva_dfm_1, sigmoid_table_861_3_sva_dfm_1, sigmoid_table_862_3_sva_dfm_1,
          sigmoid_table_863_3_sva_dfm_1, sigmoid_table_864_3_sva_dfm_1, sigmoid_table_865_3_sva_dfm_1,
          sigmoid_table_866_3_sva_dfm_1, sigmoid_table_867_2_sva_dfm_1, sigmoid_table_868_2_sva_dfm_1,
          sigmoid_table_869_2_sva_dfm_1, sigmoid_table_870_2_sva_dfm_1, sigmoid_table_871_2_sva_dfm_1,
          sigmoid_table_872_2_sva_dfm_1, sigmoid_table_873_2_sva_dfm_1, sigmoid_table_874_2_sva_dfm_1,
          sigmoid_table_875_2_sva_dfm_1, sigmoid_table_876_2_sva_dfm_1, sigmoid_table_877_2_sva_dfm_1,
          sigmoid_table_878_2_sva_dfm_1, sigmoid_table_879_2_sva_dfm_1, sigmoid_table_880_2_sva_dfm_1,
          sigmoid_table_881_2_sva_dfm_1, sigmoid_table_882_2_sva_dfm_1, sigmoid_table_883_2_sva_dfm_1,
          sigmoid_table_884_2_sva_dfm_1, sigmoid_table_885_2_sva_dfm_1, sigmoid_table_886_2_sva_dfm_1,
          sigmoid_table_887_2_sva_dfm_1, sigmoid_table_888_2_sva_dfm_1, sigmoid_table_889_2_sva_dfm_1,
          sigmoid_table_890_2_sva_dfm_1, sigmoid_table_891_2_sva_dfm_1, sigmoid_table_892_2_sva_dfm_1,
          sigmoid_table_893_2_sva_dfm_1, sigmoid_table_894_2_sva_dfm_1, sigmoid_table_895_2_sva_dfm_1,
          sigmoid_table_896_2_sva_dfm_1, sigmoid_table_897_2_sva_dfm_1, sigmoid_table_898_2_sva_dfm_1,
          sigmoid_table_899_2_sva_dfm_1, sigmoid_table_900_2_sva_dfm_1, sigmoid_table_901_2_sva_dfm_1,
          sigmoid_table_902_2_sva_dfm_1, sigmoid_table_903_2_sva_dfm_1, sigmoid_table_904_2_sva_dfm_1,
          sigmoid_table_905_2_sva_dfm_1, sigmoid_table_906_2_sva_dfm_1, sigmoid_table_907_2_sva_dfm_1,
          sigmoid_table_908_2_sva_dfm_1, sigmoid_table_909_2_sva_dfm_1, sigmoid_table_910_2_sva_dfm_1,
          sigmoid_table_911_1_sva_dfm_1, sigmoid_table_912_1_sva_dfm_1, sigmoid_table_913_1_sva_dfm_1,
          sigmoid_table_914_1_sva_dfm_1, sigmoid_table_915_1_sva_dfm_1, sigmoid_table_916_1_sva_dfm_1,
          sigmoid_table_917_1_sva_dfm_1, sigmoid_table_918_1_sva_dfm_1, sigmoid_table_919_1_sva_dfm_1,
          sigmoid_table_920_1_sva_dfm_1, sigmoid_table_921_1_sva_dfm_1, sigmoid_table_922_1_sva_dfm_1,
          sigmoid_table_923_1_sva_dfm_1, sigmoid_table_924_1_sva_dfm_1, sigmoid_table_925_1_sva_dfm_1,
          sigmoid_table_926_1_sva_dfm_1, sigmoid_table_927_1_sva_dfm_1, sigmoid_table_928_1_sva_dfm_1,
          sigmoid_table_929_1_sva_dfm_1, sigmoid_table_930_1_sva_dfm_1, sigmoid_table_931_1_sva_dfm_1,
          sigmoid_table_932_1_sva_dfm_1, sigmoid_table_933_1_sva_dfm_1, sigmoid_table_934_1_sva_dfm_1,
          sigmoid_table_935_1_sva_dfm_1, sigmoid_table_936_1_sva_dfm_1, sigmoid_table_937_1_sva_dfm_1,
          sigmoid_table_938_1_sva_dfm_1, sigmoid_table_939_1_sva_dfm_1, sigmoid_table_940_1_sva_dfm_1,
          sigmoid_table_941_1_sva_dfm_1, sigmoid_table_942_1_sva_dfm_1, sigmoid_table_943_1_sva_dfm_1,
          sigmoid_table_944_1_sva_dfm_1, sigmoid_table_945_1_sva_dfm_1, sigmoid_table_946_1_sva_dfm_1,
          sigmoid_table_947_1_sva_dfm_1, sigmoid_table_948_1_sva_dfm_1, sigmoid_table_949_1_sva_dfm_1,
          sigmoid_table_950_1_sva_dfm_1, sigmoid_table_951_1_sva_dfm_1, sigmoid_table_952_1_sva_dfm_1,
          sigmoid_table_953_1_sva_dfm_1, sigmoid_table_954_1_sva_dfm_1, sigmoid_table_955_0_sva_dfm_1,
          sigmoid_table_956_0_sva_dfm_1, sigmoid_table_957_0_sva_dfm_1, sigmoid_table_958_0_sva_dfm_1,
          sigmoid_table_959_0_sva_dfm_1, sigmoid_table_960_0_sva_dfm_1, sigmoid_table_961_0_sva_dfm_1,
          sigmoid_table_962_0_sva_dfm_1, sigmoid_table_963_0_sva_dfm_1, sigmoid_table_964_0_sva_dfm_1,
          sigmoid_table_965_0_sva_dfm_1, sigmoid_table_966_0_sva_dfm_1, sigmoid_table_967_0_sva_dfm_1,
          sigmoid_table_968_0_sva_dfm_1, sigmoid_table_969_0_sva_dfm_1, sigmoid_table_970_0_sva_dfm_1,
          sigmoid_table_971_0_sva_dfm_1, sigmoid_table_972_0_sva_dfm_1, sigmoid_table_973_0_sva_dfm_1,
          sigmoid_table_974_0_sva_dfm_1, sigmoid_table_975_0_sva_dfm_1, sigmoid_table_976_0_sva_dfm_1,
          sigmoid_table_977_0_sva_dfm_1, sigmoid_table_978_0_sva_dfm_1, sigmoid_table_979_0_sva_dfm_1,
          sigmoid_table_980_0_sva_dfm_1, sigmoid_table_981_0_sva_dfm_1, sigmoid_table_982_0_sva_dfm_1,
          sigmoid_table_983_0_sva_dfm_1, sigmoid_table_984_0_sva_dfm_1, sigmoid_table_985_0_sva_dfm_1,
          sigmoid_table_986_0_sva_dfm_1, sigmoid_table_987_0_sva_dfm_1, sigmoid_table_988_0_sva_dfm_1,
          sigmoid_table_989_0_sva_dfm_1, sigmoid_table_990_0_sva_dfm_1, sigmoid_table_991_0_sva_dfm_1,
          sigmoid_table_992_0_sva_dfm_1, sigmoid_table_993_0_sva_dfm_1, sigmoid_table_994_0_sva_dfm_1,
          sigmoid_table_995_0_sva_dfm_1, sigmoid_table_996_0_sva_dfm_1, sigmoid_table_997_0_sva_dfm_1,
          sigmoid_table_998_0_sva_dfm_1, sigmoid_table_999_0_sva_dfm_1, sigmoid_table_1000_0_sva_dfm_1,
          sigmoid_table_1001_0_sva_dfm_1, sigmoid_table_1002_0_sva_dfm_1, sigmoid_table_1003_0_sva_dfm_1,
          sigmoid_table_1004_0_sva_dfm_1, sigmoid_table_1005_0_sva_dfm_1, sigmoid_table_1006_0_sva_dfm_1,
          sigmoid_table_1007_0_sva_dfm_1, sigmoid_table_1008_0_sva_dfm_1, sigmoid_table_1009_0_sva_dfm_1,
          sigmoid_table_1010_0_sva_dfm_1, sigmoid_table_1011_0_sva_dfm_1, sigmoid_table_1012_0_sva_dfm_1,
          sigmoid_table_1013_0_sva_dfm_1, sigmoid_table_1014_0_sva_dfm_1, sigmoid_table_1015_0_sva_dfm_1,
          sigmoid_table_1016_0_sva_dfm_1, sigmoid_table_1017_0_sva_dfm_1, sigmoid_table_1018_0_sva_dfm_1,
          sigmoid_table_1019_0_sva_dfm_1, sigmoid_table_1020_0_sva_dfm_1, sigmoid_table_1021_0_sva_dfm_1,
          sigmoid_table_1022_0_sva_dfm_1, sigmoid_table_1023_0_sva_dfm_1, {for_for_or_1_itm
          , for_for_or_itm});
      res_rsci_d_2 <= MUX_s_1_1024_2(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_158_2_sva_dfm_1, sigmoid_table_159_2_sva_dfm_1,
          sigmoid_table_160_2_sva_dfm_1, sigmoid_table_161_2_sva_dfm_1, sigmoid_table_162_2_sva_dfm_1,
          sigmoid_table_163_2_sva_dfm_1, sigmoid_table_164_2_sva_dfm_1, sigmoid_table_165_2_sva_dfm_1,
          sigmoid_table_166_2_sva_dfm_1, sigmoid_table_167_2_sva_dfm_1, sigmoid_table_168_2_sva_dfm_1,
          sigmoid_table_169_2_sva_dfm_1, sigmoid_table_170_2_sva_dfm_1, sigmoid_table_171_2_sva_dfm_1,
          sigmoid_table_172_2_sva_dfm_1, sigmoid_table_173_2_sva_dfm_1, sigmoid_table_174_2_sva_dfm_1,
          sigmoid_table_175_2_sva_dfm_1, sigmoid_table_176_2_sva_dfm_1, sigmoid_table_177_2_sva_dfm_1,
          sigmoid_table_178_2_sva_dfm_1, sigmoid_table_179_2_sva_dfm_1, sigmoid_table_180_2_sva_dfm_1,
          sigmoid_table_181_2_sva_dfm_1, sigmoid_table_182_2_sva_dfm_1, sigmoid_table_183_2_sva_dfm_1,
          sigmoid_table_184_1_sva_dfm_1, sigmoid_table_185_1_sva_dfm_1, sigmoid_table_186_1_sva_dfm_1,
          sigmoid_table_187_1_sva_dfm_1, sigmoid_table_188_1_sva_dfm_1, sigmoid_table_189_1_sva_dfm_1,
          sigmoid_table_190_1_sva_dfm_1, sigmoid_table_191_1_sva_dfm_1, sigmoid_table_192_1_sva_dfm_1,
          sigmoid_table_193_1_sva_dfm_1, sigmoid_table_194_0_sva_dfm_1, sigmoid_table_195_0_sva_dfm_1,
          sigmoid_table_196_0_sva_dfm_1, sigmoid_table_197_0_sva_dfm_1, sigmoid_table_198_0_sva_dfm_1,
          sigmoid_table_199_0_sva_dfm_1, sigmoid_table_200_0_sva_dfm_1, sigmoid_table_201_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, sigmoid_table_229_2_sva_dfm_1, sigmoid_table_230_2_sva_dfm_1,
          sigmoid_table_231_2_sva_dfm_1, sigmoid_table_232_2_sva_dfm_1, sigmoid_table_233_2_sva_dfm_1,
          sigmoid_table_234_2_sva_dfm_1, sigmoid_table_235_2_sva_dfm_1, sigmoid_table_236_2_sva_dfm_1,
          sigmoid_table_237_2_sva_dfm_1, sigmoid_table_238_2_sva_dfm_1, sigmoid_table_239_1_sva_dfm_1,
          sigmoid_table_240_1_sva_dfm_1, sigmoid_table_241_1_sva_dfm_1, sigmoid_table_242_1_sva_dfm_1,
          sigmoid_table_243_0_sva_dfm_1, sigmoid_table_244_0_sva_dfm_1, sigmoid_table_245_0_sva_dfm_1,
          sigmoid_table_246_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_262_2_sva_dfm_1,
          sigmoid_table_263_2_sva_dfm_1, sigmoid_table_264_2_sva_dfm_1, sigmoid_table_265_2_sva_dfm_1,
          sigmoid_table_266_2_sva_dfm_1, sigmoid_table_267_2_sva_dfm_1, sigmoid_table_268_1_sva_dfm_1,
          sigmoid_table_269_1_sva_dfm_1, sigmoid_table_270_1_sva_dfm_1, sigmoid_table_271_0_sva_dfm_1,
          sigmoid_table_272_0_sva_dfm_1, sigmoid_table_273_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_284_2_sva_dfm_1,
          sigmoid_table_285_2_sva_dfm_1, sigmoid_table_286_2_sva_dfm_1, sigmoid_table_287_2_sva_dfm_1,
          sigmoid_table_288_1_sva_dfm_1, sigmoid_table_289_1_sva_dfm_1, sigmoid_table_290_1_sva_dfm_1,
          sigmoid_table_291_0_sva_dfm_1, sigmoid_table_292_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_301_2_sva_dfm_1, sigmoid_table_302_2_sva_dfm_1,
          sigmoid_table_303_2_sva_dfm_1, sigmoid_table_304_1_sva_dfm_1, sigmoid_table_305_1_sva_dfm_1,
          sigmoid_table_306_0_sva_dfm_1, sigmoid_table_307_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_314_2_sva_dfm_1, sigmoid_table_315_2_sva_dfm_1,
          sigmoid_table_316_2_sva_dfm_1, sigmoid_table_317_1_sva_dfm_1, sigmoid_table_318_0_sva_dfm_1,
          sigmoid_table_319_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_325_2_sva_dfm_1,
          sigmoid_table_326_2_sva_dfm_1, sigmoid_table_327_2_sva_dfm_1, sigmoid_table_328_1_sva_dfm_1,
          sigmoid_table_329_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_335_2_sva_dfm_1,
          sigmoid_table_336_2_sva_dfm_1, sigmoid_table_337_1_sva_dfm_1, sigmoid_table_338_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_343_2_sva_dfm_1, sigmoid_table_344_2_sva_dfm_1,
          sigmoid_table_345_1_sva_dfm_1, sigmoid_table_346_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_351_2_sva_dfm_1, sigmoid_table_352_2_sva_dfm_1,
          sigmoid_table_353_1_sva_dfm_1, sigmoid_table_354_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, sigmoid_table_358_2_sva_dfm_1, sigmoid_table_359_2_sva_dfm_1, sigmoid_table_360_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, sigmoid_table_364_2_sva_dfm_1, sigmoid_table_365_2_sva_dfm_1,
          sigmoid_table_366_1_sva_dfm_1, 1'b0, 1'b0, 1'b0, sigmoid_table_370_2_sva_dfm_1,
          sigmoid_table_371_2_sva_dfm_1, sigmoid_table_372_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, sigmoid_table_376_2_sva_dfm_1, sigmoid_table_377_1_sva_dfm_1, 1'b0,
          1'b0, 1'b0, sigmoid_table_381_2_sva_dfm_1, sigmoid_table_382_1_sva_dfm_1,
          1'b0, 1'b0, 1'b0, sigmoid_table_386_2_sva_dfm_1, sigmoid_table_387_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_390_2_sva_dfm_1, sigmoid_table_391_1_sva_dfm_1,
          1'b0, 1'b0, 1'b0, sigmoid_table_395_2_sva_dfm_1, sigmoid_table_396_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_399_2_sva_dfm_1, sigmoid_table_400_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_403_2_sva_dfm_1, sigmoid_table_404_0_sva_dfm_1,
          1'b0, sigmoid_table_406_2_sva_dfm_1, sigmoid_table_407_1_sva_dfm_1, 1'b0,
          1'b0, sigmoid_table_410_2_sva_dfm_1, sigmoid_table_411_0_sva_dfm_1, 1'b0,
          1'b0, sigmoid_table_414_1_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_417_2_sva_dfm_1,
          sigmoid_table_418_0_sva_dfm_1, 1'b0, sigmoid_table_420_2_sva_dfm_1, sigmoid_table_421_0_sva_dfm_1,
          1'b0, sigmoid_table_423_2_sva_dfm_1, sigmoid_table_424_1_sva_dfm_1, 1'b0,
          1'b0, sigmoid_table_427_1_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_430_1_sva_dfm_1,
          1'b0, sigmoid_table_432_2_sva_dfm_1, sigmoid_table_433_1_sva_dfm_1, 1'b0,
          sigmoid_table_435_2_sva_dfm_1, sigmoid_table_436_0_sva_dfm_1, 1'b0, sigmoid_table_438_2_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_441_2_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_444_1_sva_dfm_1,
          1'b0, sigmoid_table_446_2_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_449_1_sva_dfm_1,
          1'b0, sigmoid_table_451_2_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_454_1_sva_dfm_1,
          1'b0, sigmoid_table_456_2_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_459_0_sva_dfm_1,
          1'b0, sigmoid_table_461_1_sva_dfm_1, 1'b0, sigmoid_table_463_2_sva_dfm_1,
          1'b0, sigmoid_table_465_2_sva_dfm_1, sigmoid_table_466_0_sva_dfm_1, 1'b0,
          sigmoid_table_468_1_sva_dfm_1, 1'b0, sigmoid_table_470_2_sva_dfm_1, 1'b0,
          sigmoid_table_472_2_sva_dfm_1, 1'b0, sigmoid_table_474_2_sva_dfm_1, sigmoid_table_475_0_sva_dfm_1,
          1'b0, sigmoid_table_477_0_sva_dfm_1, 1'b0, sigmoid_table_479_1_sva_dfm_1,
          1'b0, sigmoid_table_481_1_sva_dfm_1, 1'b0, sigmoid_table_483_2_sva_dfm_1,
          1'b0, sigmoid_table_485_2_sva_dfm_1, 1'b0, sigmoid_table_487_2_sva_dfm_1,
          1'b0, sigmoid_table_489_2_sva_dfm_1, 1'b0, sigmoid_table_491_2_sva_dfm_1,
          1'b0, sigmoid_table_493_2_sva_dfm_1, 1'b0, sigmoid_table_495_2_sva_dfm_1,
          1'b0, sigmoid_table_497_2_sva_dfm_1, 1'b0, sigmoid_table_499_2_sva_dfm_1,
          1'b0, sigmoid_table_501_2_sva_dfm_1, 1'b0, sigmoid_table_503_2_sva_dfm_1,
          1'b0, sigmoid_table_505_2_sva_dfm_1, 1'b0, sigmoid_table_507_2_sva_dfm_1,
          1'b0, sigmoid_table_509_2_sva_dfm_1, 1'b0, sigmoid_table_511_2_sva_dfm_1,
          1'b0, sigmoid_table_513_2_sva_dfm_1, 1'b0, sigmoid_table_515_2_sva_dfm_1,
          sigmoid_table_516_0_sva_dfm_1, 1'b0, sigmoid_table_518_0_sva_dfm_1, 1'b0,
          sigmoid_table_520_0_sva_dfm_1, 1'b0, sigmoid_table_522_0_sva_dfm_1, 1'b0,
          sigmoid_table_524_0_sva_dfm_1, 1'b0, sigmoid_table_526_0_sva_dfm_1, 1'b0,
          sigmoid_table_528_0_sva_dfm_1, 1'b0, sigmoid_table_530_0_sva_dfm_1, 1'b0,
          sigmoid_table_532_0_sva_dfm_1, 1'b0, sigmoid_table_534_0_sva_dfm_1, 1'b0,
          sigmoid_table_536_1_sva_dfm_1, 1'b0, sigmoid_table_538_1_sva_dfm_1, 1'b0,
          sigmoid_table_540_1_sva_dfm_1, 1'b0, sigmoid_table_542_2_sva_dfm_1, 1'b0,
          sigmoid_table_544_2_sva_dfm_1, 1'b0, sigmoid_table_546_2_sva_dfm_1, 1'b0,
          sigmoid_table_548_2_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_551_0_sva_dfm_1,
          1'b0, sigmoid_table_553_1_sva_dfm_1, 1'b0, sigmoid_table_555_2_sva_dfm_1,
          1'b0, sigmoid_table_557_2_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_560_0_sva_dfm_1,
          1'b0, sigmoid_table_562_1_sva_dfm_1, 1'b0, sigmoid_table_564_2_sva_dfm_1,
          1'b0, sigmoid_table_566_2_sva_dfm_1, sigmoid_table_567_0_sva_dfm_1, 1'b0,
          sigmoid_table_569_1_sva_dfm_1, 1'b0, sigmoid_table_571_2_sva_dfm_1, sigmoid_table_572_0_sva_dfm_1,
          1'b0, sigmoid_table_574_1_sva_dfm_1, 1'b0, sigmoid_table_576_2_sva_dfm_1,
          sigmoid_table_577_0_sva_dfm_1, 1'b0, sigmoid_table_579_2_sva_dfm_1, 1'b0,
          sigmoid_table_581_2_sva_dfm_1, sigmoid_table_582_0_sva_dfm_1, 1'b0, sigmoid_table_584_2_sva_dfm_1,
          sigmoid_table_585_0_sva_dfm_1, 1'b0, sigmoid_table_587_2_sva_dfm_1, 1'b0,
          1'b0, sigmoid_table_590_1_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_593_1_sva_dfm_1,
          1'b0, sigmoid_table_595_2_sva_dfm_1, sigmoid_table_596_1_sva_dfm_1, 1'b0,
          sigmoid_table_598_2_sva_dfm_1, sigmoid_table_599_1_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_602_1_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_605_2_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_608_2_sva_dfm_1, sigmoid_table_609_0_sva_dfm_1,
          1'b0, sigmoid_table_611_2_sva_dfm_1, sigmoid_table_612_1_sva_dfm_1, 1'b0,
          1'b0, sigmoid_table_615_2_sva_dfm_1, sigmoid_table_616_0_sva_dfm_1, 1'b0,
          1'b0, sigmoid_table_619_1_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_622_2_sva_dfm_1,
          sigmoid_table_623_1_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_626_2_sva_dfm_1,
          sigmoid_table_627_1_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_630_2_sva_dfm_1,
          sigmoid_table_631_2_sva_dfm_1, sigmoid_table_632_0_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_635_2_sva_dfm_1, sigmoid_table_636_0_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_639_2_sva_dfm_1, sigmoid_table_640_2_sva_dfm_1, sigmoid_table_641_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_644_2_sva_dfm_1, sigmoid_table_645_1_sva_dfm_1,
          sigmoid_table_646_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_649_2_sva_dfm_1,
          sigmoid_table_650_2_sva_dfm_1, sigmoid_table_651_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, sigmoid_table_655_2_sva_dfm_1, sigmoid_table_656_1_sva_dfm_1, sigmoid_table_657_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, sigmoid_table_661_2_sva_dfm_1, sigmoid_table_662_1_sva_dfm_1,
          sigmoid_table_663_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, sigmoid_table_667_2_sva_dfm_1,
          sigmoid_table_668_2_sva_dfm_1, sigmoid_table_669_1_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_674_2_sva_dfm_1, sigmoid_table_675_2_sva_dfm_1,
          sigmoid_table_676_1_sva_dfm_1, sigmoid_table_677_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_682_2_sva_dfm_1, sigmoid_table_683_2_sva_dfm_1,
          sigmoid_table_684_1_sva_dfm_1, sigmoid_table_685_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_690_2_sva_dfm_1, sigmoid_table_691_2_sva_dfm_1,
          sigmoid_table_692_2_sva_dfm_1, sigmoid_table_693_1_sva_dfm_1, sigmoid_table_694_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_700_2_sva_dfm_1, sigmoid_table_701_2_sva_dfm_1,
          sigmoid_table_702_2_sva_dfm_1, sigmoid_table_703_1_sva_dfm_1, sigmoid_table_704_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_711_2_sva_dfm_1, sigmoid_table_712_2_sva_dfm_1,
          sigmoid_table_713_2_sva_dfm_1, sigmoid_table_714_1_sva_dfm_1, sigmoid_table_715_1_sva_dfm_1,
          sigmoid_table_716_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          sigmoid_table_724_2_sva_dfm_1, sigmoid_table_725_2_sva_dfm_1, sigmoid_table_726_2_sva_dfm_1,
          sigmoid_table_727_2_sva_dfm_1, sigmoid_table_728_1_sva_dfm_1, sigmoid_table_729_1_sva_dfm_1,
          sigmoid_table_730_0_sva_dfm_1, sigmoid_table_731_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_741_2_sva_dfm_1,
          sigmoid_table_742_2_sva_dfm_1, sigmoid_table_743_2_sva_dfm_1, sigmoid_table_744_2_sva_dfm_1,
          sigmoid_table_745_2_sva_dfm_1, sigmoid_table_746_1_sva_dfm_1, sigmoid_table_747_1_sva_dfm_1,
          sigmoid_table_748_0_sva_dfm_1, sigmoid_table_749_0_sva_dfm_1, sigmoid_table_750_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          sigmoid_table_763_2_sva_dfm_1, sigmoid_table_764_2_sva_dfm_1, sigmoid_table_765_2_sva_dfm_1,
          sigmoid_table_766_2_sva_dfm_1, sigmoid_table_767_2_sva_dfm_1, sigmoid_table_768_2_sva_dfm_1,
          sigmoid_table_769_2_sva_dfm_1, sigmoid_table_770_1_sva_dfm_1, sigmoid_table_771_1_sva_dfm_1,
          sigmoid_table_772_1_sva_dfm_1, sigmoid_table_773_1_sva_dfm_1, sigmoid_table_774_0_sva_dfm_1,
          sigmoid_table_775_0_sva_dfm_1, sigmoid_table_776_0_sva_dfm_1, sigmoid_table_777_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_796_2_sva_dfm_1, sigmoid_table_797_2_sva_dfm_1,
          sigmoid_table_798_2_sva_dfm_1, sigmoid_table_799_2_sva_dfm_1, sigmoid_table_800_2_sva_dfm_1,
          sigmoid_table_801_2_sva_dfm_1, sigmoid_table_802_2_sva_dfm_1, sigmoid_table_803_2_sva_dfm_1,
          sigmoid_table_804_2_sva_dfm_1, sigmoid_table_805_2_sva_dfm_1, sigmoid_table_806_2_sva_dfm_1,
          sigmoid_table_807_2_sva_dfm_1, sigmoid_table_808_1_sva_dfm_1, sigmoid_table_809_1_sva_dfm_1,
          sigmoid_table_810_1_sva_dfm_1, sigmoid_table_811_1_sva_dfm_1, sigmoid_table_812_1_sva_dfm_1,
          sigmoid_table_813_1_sva_dfm_1, sigmoid_table_814_1_sva_dfm_1, sigmoid_table_815_0_sva_dfm_1,
          sigmoid_table_816_0_sva_dfm_1, sigmoid_table_817_0_sva_dfm_1, sigmoid_table_818_0_sva_dfm_1,
          sigmoid_table_819_0_sva_dfm_1, sigmoid_table_820_0_sva_dfm_1, sigmoid_table_821_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_867_2_sva_dfm_1,
          sigmoid_table_868_2_sva_dfm_1, sigmoid_table_869_2_sva_dfm_1, sigmoid_table_870_2_sva_dfm_1,
          sigmoid_table_871_2_sva_dfm_1, sigmoid_table_872_2_sva_dfm_1, sigmoid_table_873_2_sva_dfm_1,
          sigmoid_table_874_2_sva_dfm_1, sigmoid_table_875_2_sva_dfm_1, sigmoid_table_876_2_sva_dfm_1,
          sigmoid_table_877_2_sva_dfm_1, sigmoid_table_878_2_sva_dfm_1, sigmoid_table_879_2_sva_dfm_1,
          sigmoid_table_880_2_sva_dfm_1, sigmoid_table_881_2_sva_dfm_1, sigmoid_table_882_2_sva_dfm_1,
          sigmoid_table_883_2_sva_dfm_1, sigmoid_table_884_2_sva_dfm_1, sigmoid_table_885_2_sva_dfm_1,
          sigmoid_table_886_2_sva_dfm_1, sigmoid_table_887_2_sva_dfm_1, sigmoid_table_888_2_sva_dfm_1,
          sigmoid_table_889_2_sva_dfm_1, sigmoid_table_890_2_sva_dfm_1, sigmoid_table_891_2_sva_dfm_1,
          sigmoid_table_892_2_sva_dfm_1, sigmoid_table_893_2_sva_dfm_1, sigmoid_table_894_2_sva_dfm_1,
          sigmoid_table_895_2_sva_dfm_1, sigmoid_table_896_2_sva_dfm_1, sigmoid_table_897_2_sva_dfm_1,
          sigmoid_table_898_2_sva_dfm_1, sigmoid_table_899_2_sva_dfm_1, sigmoid_table_900_2_sva_dfm_1,
          sigmoid_table_901_2_sva_dfm_1, sigmoid_table_902_2_sva_dfm_1, sigmoid_table_903_2_sva_dfm_1,
          sigmoid_table_904_2_sva_dfm_1, sigmoid_table_905_2_sva_dfm_1, sigmoid_table_906_2_sva_dfm_1,
          sigmoid_table_907_2_sva_dfm_1, sigmoid_table_908_2_sva_dfm_1, sigmoid_table_909_2_sva_dfm_1,
          sigmoid_table_910_2_sva_dfm_1, sigmoid_table_911_1_sva_dfm_1, sigmoid_table_912_1_sva_dfm_1,
          sigmoid_table_913_1_sva_dfm_1, sigmoid_table_914_1_sva_dfm_1, sigmoid_table_915_1_sva_dfm_1,
          sigmoid_table_916_1_sva_dfm_1, sigmoid_table_917_1_sva_dfm_1, sigmoid_table_918_1_sva_dfm_1,
          sigmoid_table_919_1_sva_dfm_1, sigmoid_table_920_1_sva_dfm_1, sigmoid_table_921_1_sva_dfm_1,
          sigmoid_table_922_1_sva_dfm_1, sigmoid_table_923_1_sva_dfm_1, sigmoid_table_924_1_sva_dfm_1,
          sigmoid_table_925_1_sva_dfm_1, sigmoid_table_926_1_sva_dfm_1, sigmoid_table_927_1_sva_dfm_1,
          sigmoid_table_928_1_sva_dfm_1, sigmoid_table_929_1_sva_dfm_1, sigmoid_table_930_1_sva_dfm_1,
          sigmoid_table_931_1_sva_dfm_1, sigmoid_table_932_1_sva_dfm_1, sigmoid_table_933_1_sva_dfm_1,
          sigmoid_table_934_1_sva_dfm_1, sigmoid_table_935_1_sva_dfm_1, sigmoid_table_936_1_sva_dfm_1,
          sigmoid_table_937_1_sva_dfm_1, sigmoid_table_938_1_sva_dfm_1, sigmoid_table_939_1_sva_dfm_1,
          sigmoid_table_940_1_sva_dfm_1, sigmoid_table_941_1_sva_dfm_1, sigmoid_table_942_1_sva_dfm_1,
          sigmoid_table_943_1_sva_dfm_1, sigmoid_table_944_1_sva_dfm_1, sigmoid_table_945_1_sva_dfm_1,
          sigmoid_table_946_1_sva_dfm_1, sigmoid_table_947_1_sva_dfm_1, sigmoid_table_948_1_sva_dfm_1,
          sigmoid_table_949_1_sva_dfm_1, sigmoid_table_950_1_sva_dfm_1, sigmoid_table_951_1_sva_dfm_1,
          sigmoid_table_952_1_sva_dfm_1, sigmoid_table_953_1_sva_dfm_1, sigmoid_table_954_1_sva_dfm_1,
          sigmoid_table_955_0_sva_dfm_1, sigmoid_table_956_0_sva_dfm_1, sigmoid_table_957_0_sva_dfm_1,
          sigmoid_table_958_0_sva_dfm_1, sigmoid_table_959_0_sva_dfm_1, sigmoid_table_960_0_sva_dfm_1,
          sigmoid_table_961_0_sva_dfm_1, sigmoid_table_962_0_sva_dfm_1, sigmoid_table_963_0_sva_dfm_1,
          sigmoid_table_964_0_sva_dfm_1, sigmoid_table_965_0_sva_dfm_1, sigmoid_table_966_0_sva_dfm_1,
          sigmoid_table_967_0_sva_dfm_1, sigmoid_table_968_0_sva_dfm_1, sigmoid_table_969_0_sva_dfm_1,
          sigmoid_table_970_0_sva_dfm_1, sigmoid_table_971_0_sva_dfm_1, sigmoid_table_972_0_sva_dfm_1,
          sigmoid_table_973_0_sva_dfm_1, sigmoid_table_974_0_sva_dfm_1, sigmoid_table_975_0_sva_dfm_1,
          sigmoid_table_976_0_sva_dfm_1, sigmoid_table_977_0_sva_dfm_1, sigmoid_table_978_0_sva_dfm_1,
          sigmoid_table_979_0_sva_dfm_1, sigmoid_table_980_0_sva_dfm_1, sigmoid_table_981_0_sva_dfm_1,
          sigmoid_table_982_0_sva_dfm_1, sigmoid_table_983_0_sva_dfm_1, sigmoid_table_984_0_sva_dfm_1,
          sigmoid_table_985_0_sva_dfm_1, sigmoid_table_986_0_sva_dfm_1, sigmoid_table_987_0_sva_dfm_1,
          sigmoid_table_988_0_sva_dfm_1, sigmoid_table_989_0_sva_dfm_1, sigmoid_table_990_0_sva_dfm_1,
          sigmoid_table_991_0_sva_dfm_1, sigmoid_table_992_0_sva_dfm_1, sigmoid_table_993_0_sva_dfm_1,
          sigmoid_table_994_0_sva_dfm_1, sigmoid_table_995_0_sva_dfm_1, sigmoid_table_996_0_sva_dfm_1,
          sigmoid_table_997_0_sva_dfm_1, sigmoid_table_998_0_sva_dfm_1, sigmoid_table_999_0_sva_dfm_1,
          sigmoid_table_1000_0_sva_dfm_1, sigmoid_table_1001_0_sva_dfm_1, sigmoid_table_1002_0_sva_dfm_1,
          sigmoid_table_1003_0_sva_dfm_1, sigmoid_table_1004_0_sva_dfm_1, sigmoid_table_1005_0_sva_dfm_1,
          sigmoid_table_1006_0_sva_dfm_1, sigmoid_table_1007_0_sva_dfm_1, sigmoid_table_1008_0_sva_dfm_1,
          sigmoid_table_1009_0_sva_dfm_1, sigmoid_table_1010_0_sva_dfm_1, sigmoid_table_1011_0_sva_dfm_1,
          sigmoid_table_1012_0_sva_dfm_1, sigmoid_table_1013_0_sva_dfm_1, sigmoid_table_1014_0_sva_dfm_1,
          sigmoid_table_1015_0_sva_dfm_1, sigmoid_table_1016_0_sva_dfm_1, sigmoid_table_1017_0_sva_dfm_1,
          sigmoid_table_1018_0_sva_dfm_1, sigmoid_table_1019_0_sva_dfm_1, sigmoid_table_1020_0_sva_dfm_1,
          sigmoid_table_1021_0_sva_dfm_1, sigmoid_table_1022_0_sva_dfm_1, sigmoid_table_1023_0_sva_dfm_1,
          {for_for_or_1_itm , for_for_or_itm});
      res_rsci_d_7 <= MUX_s_1_1024_2(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_388_7_sva_dfm_1,
          sigmoid_table_389_7_sva_dfm_1, sigmoid_table_390_7_sva_dfm_1, sigmoid_table_391_7_sva_dfm_1,
          sigmoid_table_392_7_sva_dfm_1, sigmoid_table_393_7_sva_dfm_1, sigmoid_table_394_7_sva_dfm_1,
          sigmoid_table_395_7_sva_dfm_1, sigmoid_table_396_7_sva_dfm_1, sigmoid_table_397_7_sva_dfm_1,
          sigmoid_table_398_7_sva_dfm_1, sigmoid_table_399_7_sva_dfm_1, sigmoid_table_400_7_sva_dfm_1,
          sigmoid_table_401_7_sva_dfm_1, sigmoid_table_402_7_sva_dfm_1, sigmoid_table_403_7_sva_dfm_1,
          sigmoid_table_404_7_sva_dfm_1, sigmoid_table_405_7_sva_dfm_1, sigmoid_table_406_7_sva_dfm_1,
          sigmoid_table_407_7_sva_dfm_1, sigmoid_table_408_7_sva_dfm_1, sigmoid_table_409_7_sva_dfm_1,
          sigmoid_table_410_7_sva_dfm_1, sigmoid_table_411_7_sva_dfm_1, sigmoid_table_412_7_sva_dfm_1,
          sigmoid_table_413_7_sva_dfm_1, sigmoid_table_414_7_sva_dfm_1, sigmoid_table_415_7_sva_dfm_1,
          sigmoid_table_416_7_sva_dfm_1, sigmoid_table_417_7_sva_dfm_1, sigmoid_table_418_7_sva_dfm_1,
          sigmoid_table_419_6_sva_dfm_1, sigmoid_table_420_6_sva_dfm_1, sigmoid_table_421_6_sva_dfm_1,
          sigmoid_table_422_6_sva_dfm_1, sigmoid_table_423_6_sva_dfm_1, sigmoid_table_424_6_sva_dfm_1,
          sigmoid_table_425_6_sva_dfm_1, sigmoid_table_426_6_sva_dfm_1, sigmoid_table_427_6_sva_dfm_1,
          sigmoid_table_428_6_sva_dfm_1, sigmoid_table_429_6_sva_dfm_1, sigmoid_table_430_6_sva_dfm_1,
          sigmoid_table_431_5_sva_dfm_1, sigmoid_table_432_5_sva_dfm_1, sigmoid_table_433_5_sva_dfm_1,
          sigmoid_table_434_5_sva_dfm_1, sigmoid_table_435_5_sva_dfm_1, sigmoid_table_436_5_sva_dfm_1,
          sigmoid_table_437_4_sva_dfm_1, sigmoid_table_438_4_sva_dfm_1, sigmoid_table_439_3_sva_dfm_1,
          sigmoid_table_440_3_sva_dfm_1, sigmoid_table_441_2_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          sigmoid_table_480_7_sva_dfm_1, sigmoid_table_481_7_sva_dfm_1, sigmoid_table_482_7_sva_dfm_1,
          sigmoid_table_483_7_sva_dfm_1, sigmoid_table_484_7_sva_dfm_1, sigmoid_table_485_7_sva_dfm_1,
          sigmoid_table_486_7_sva_dfm_1, sigmoid_table_487_7_sva_dfm_1, sigmoid_table_488_7_sva_dfm_1,
          sigmoid_table_489_7_sva_dfm_1, sigmoid_table_490_7_sva_dfm_1, sigmoid_table_491_7_sva_dfm_1,
          sigmoid_table_492_7_sva_dfm_1, sigmoid_table_493_7_sva_dfm_1, sigmoid_table_494_7_sva_dfm_1,
          sigmoid_table_495_7_sva_dfm_1, sigmoid_table_496_6_sva_dfm_1, sigmoid_table_497_6_sva_dfm_1,
          sigmoid_table_498_6_sva_dfm_1, sigmoid_table_499_6_sva_dfm_1, sigmoid_table_500_6_sva_dfm_1,
          sigmoid_table_501_6_sva_dfm_1, sigmoid_table_502_6_sva_dfm_1, sigmoid_table_503_6_sva_dfm_1,
          sigmoid_table_504_5_sva_dfm_1, sigmoid_table_505_5_sva_dfm_1, sigmoid_table_506_5_sva_dfm_1,
          sigmoid_table_507_5_sva_dfm_1, sigmoid_table_508_4_sva_dfm_1, sigmoid_table_509_4_sva_dfm_1,
          sigmoid_table_510_3_sva_dfm_1, sigmoid_table_511_2_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_545_7_sva_dfm_1,
          sigmoid_table_546_7_sva_dfm_1, sigmoid_table_547_7_sva_dfm_1, sigmoid_table_548_7_sva_dfm_1,
          sigmoid_table_549_7_sva_dfm_1, sigmoid_table_550_7_sva_dfm_1, sigmoid_table_551_7_sva_dfm_1,
          sigmoid_table_552_7_sva_dfm_1, sigmoid_table_553_7_sva_dfm_1, sigmoid_table_554_7_sva_dfm_1,
          sigmoid_table_555_7_sva_dfm_1, sigmoid_table_556_7_sva_dfm_1, sigmoid_table_557_7_sva_dfm_1,
          sigmoid_table_558_7_sva_dfm_1, sigmoid_table_559_7_sva_dfm_1, sigmoid_table_560_7_sva_dfm_1,
          sigmoid_table_561_7_sva_dfm_1, sigmoid_table_562_7_sva_dfm_1, sigmoid_table_563_6_sva_dfm_1,
          sigmoid_table_564_6_sva_dfm_1, sigmoid_table_565_6_sva_dfm_1, sigmoid_table_566_6_sva_dfm_1,
          sigmoid_table_567_6_sva_dfm_1, sigmoid_table_568_6_sva_dfm_1, sigmoid_table_569_6_sva_dfm_1,
          sigmoid_table_570_6_sva_dfm_1, sigmoid_table_571_6_sva_dfm_1, sigmoid_table_572_6_sva_dfm_1,
          sigmoid_table_573_5_sva_dfm_1, sigmoid_table_574_5_sva_dfm_1, sigmoid_table_575_5_sva_dfm_1,
          sigmoid_table_576_5_sva_dfm_1, sigmoid_table_577_5_sva_dfm_1, sigmoid_table_578_4_sva_dfm_1,
          sigmoid_table_579_4_sva_dfm_1, sigmoid_table_580_3_sva_dfm_1, sigmoid_table_581_2_sva_dfm_1,
          sigmoid_table_582_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_637_7_sva_dfm_1,
          sigmoid_table_638_7_sva_dfm_1, sigmoid_table_639_7_sva_dfm_1, sigmoid_table_640_7_sva_dfm_1,
          sigmoid_table_641_7_sva_dfm_1, sigmoid_table_642_7_sva_dfm_1, sigmoid_table_643_7_sva_dfm_1,
          sigmoid_table_644_7_sva_dfm_1, sigmoid_table_645_7_sva_dfm_1, sigmoid_table_646_7_sva_dfm_1,
          sigmoid_table_647_7_sva_dfm_1, sigmoid_table_648_7_sva_dfm_1, sigmoid_table_649_7_sva_dfm_1,
          sigmoid_table_650_7_sva_dfm_1, sigmoid_table_651_7_sva_dfm_1, sigmoid_table_652_7_sva_dfm_1,
          sigmoid_table_653_7_sva_dfm_1, sigmoid_table_654_7_sva_dfm_1, sigmoid_table_655_7_sva_dfm_1,
          sigmoid_table_656_7_sva_dfm_1, sigmoid_table_657_7_sva_dfm_1, sigmoid_table_658_7_sva_dfm_1,
          sigmoid_table_659_7_sva_dfm_1, sigmoid_table_660_7_sva_dfm_1, sigmoid_table_661_7_sva_dfm_1,
          sigmoid_table_662_7_sva_dfm_1, sigmoid_table_663_7_sva_dfm_1, sigmoid_table_664_7_sva_dfm_1,
          sigmoid_table_665_7_sva_dfm_1, sigmoid_table_666_7_sva_dfm_1, sigmoid_table_667_7_sva_dfm_1,
          sigmoid_table_668_7_sva_dfm_1, sigmoid_table_669_7_sva_dfm_1, sigmoid_table_670_7_sva_dfm_1,
          sigmoid_table_671_7_sva_dfm_1, sigmoid_table_672_7_sva_dfm_1, sigmoid_table_673_7_sva_dfm_1,
          sigmoid_table_674_7_sva_dfm_1, sigmoid_table_675_7_sva_dfm_1, sigmoid_table_676_7_sva_dfm_1,
          sigmoid_table_677_7_sva_dfm_1, sigmoid_table_678_7_sva_dfm_1, sigmoid_table_679_7_sva_dfm_1,
          sigmoid_table_680_7_sva_dfm_1, sigmoid_table_681_7_sva_dfm_1, sigmoid_table_682_7_sva_dfm_1,
          sigmoid_table_683_7_sva_dfm_1, sigmoid_table_684_7_sva_dfm_1, sigmoid_table_685_7_sva_dfm_1,
          sigmoid_table_686_6_sva_dfm_1, sigmoid_table_687_6_sva_dfm_1, sigmoid_table_688_6_sva_dfm_1,
          sigmoid_table_689_6_sva_dfm_1, sigmoid_table_690_6_sva_dfm_1, sigmoid_table_691_6_sva_dfm_1,
          sigmoid_table_692_6_sva_dfm_1, sigmoid_table_693_6_sva_dfm_1, sigmoid_table_694_6_sva_dfm_1,
          sigmoid_table_695_6_sva_dfm_1, sigmoid_table_696_6_sva_dfm_1, sigmoid_table_697_6_sva_dfm_1,
          sigmoid_table_698_6_sva_dfm_1, sigmoid_table_699_6_sva_dfm_1, sigmoid_table_700_6_sva_dfm_1,
          sigmoid_table_701_6_sva_dfm_1, sigmoid_table_702_6_sva_dfm_1, sigmoid_table_703_6_sva_dfm_1,
          sigmoid_table_704_6_sva_dfm_1, sigmoid_table_705_6_sva_dfm_1, sigmoid_table_706_6_sva_dfm_1,
          sigmoid_table_707_6_sva_dfm_1, sigmoid_table_708_6_sva_dfm_1, sigmoid_table_709_6_sva_dfm_1,
          sigmoid_table_710_6_sva_dfm_1, sigmoid_table_711_6_sva_dfm_1, sigmoid_table_712_6_sva_dfm_1,
          sigmoid_table_713_6_sva_dfm_1, sigmoid_table_714_6_sva_dfm_1, sigmoid_table_715_6_sva_dfm_1,
          sigmoid_table_716_6_sva_dfm_1, sigmoid_table_717_6_sva_dfm_1, sigmoid_table_718_6_sva_dfm_1,
          sigmoid_table_719_6_sva_dfm_1, sigmoid_table_720_6_sva_dfm_1, sigmoid_table_721_6_sva_dfm_1,
          sigmoid_table_722_6_sva_dfm_1, sigmoid_table_723_6_sva_dfm_1, sigmoid_table_724_6_sva_dfm_1,
          sigmoid_table_725_6_sva_dfm_1, sigmoid_table_726_6_sva_dfm_1, sigmoid_table_727_6_sva_dfm_1,
          sigmoid_table_728_6_sva_dfm_1, sigmoid_table_729_6_sva_dfm_1, sigmoid_table_730_6_sva_dfm_1,
          sigmoid_table_731_6_sva_dfm_1, sigmoid_table_732_5_sva_dfm_1, sigmoid_table_733_5_sva_dfm_1,
          sigmoid_table_734_5_sva_dfm_1, sigmoid_table_735_5_sva_dfm_1, sigmoid_table_736_5_sva_dfm_1,
          sigmoid_table_737_5_sva_dfm_1, sigmoid_table_738_5_sva_dfm_1, sigmoid_table_739_5_sva_dfm_1,
          sigmoid_table_740_5_sva_dfm_1, sigmoid_table_741_5_sva_dfm_1, sigmoid_table_742_5_sva_dfm_1,
          sigmoid_table_743_5_sva_dfm_1, sigmoid_table_744_5_sva_dfm_1, sigmoid_table_745_5_sva_dfm_1,
          sigmoid_table_746_5_sva_dfm_1, sigmoid_table_747_5_sva_dfm_1, sigmoid_table_748_5_sva_dfm_1,
          sigmoid_table_749_5_sva_dfm_1, sigmoid_table_750_5_sva_dfm_1, sigmoid_table_751_5_sva_dfm_1,
          sigmoid_table_752_5_sva_dfm_1, sigmoid_table_753_5_sva_dfm_1, sigmoid_table_754_5_sva_dfm_1,
          sigmoid_table_755_5_sva_dfm_1, sigmoid_table_756_5_sva_dfm_1, sigmoid_table_757_5_sva_dfm_1,
          sigmoid_table_758_5_sva_dfm_1, sigmoid_table_759_5_sva_dfm_1, sigmoid_table_760_5_sva_dfm_1,
          sigmoid_table_761_5_sva_dfm_1, sigmoid_table_762_5_sva_dfm_1, sigmoid_table_763_5_sva_dfm_1,
          sigmoid_table_764_5_sva_dfm_1, sigmoid_table_765_5_sva_dfm_1, sigmoid_table_766_5_sva_dfm_1,
          sigmoid_table_767_5_sva_dfm_1, sigmoid_table_768_5_sva_dfm_1, sigmoid_table_769_5_sva_dfm_1,
          sigmoid_table_770_5_sva_dfm_1, sigmoid_table_771_5_sva_dfm_1, sigmoid_table_772_5_sva_dfm_1,
          sigmoid_table_773_5_sva_dfm_1, sigmoid_table_774_5_sva_dfm_1, sigmoid_table_775_5_sva_dfm_1,
          sigmoid_table_776_5_sva_dfm_1, sigmoid_table_777_5_sva_dfm_1, sigmoid_table_778_4_sva_dfm_1,
          sigmoid_table_779_4_sva_dfm_1, sigmoid_table_780_4_sva_dfm_1, sigmoid_table_781_4_sva_dfm_1,
          sigmoid_table_782_4_sva_dfm_1, sigmoid_table_783_4_sva_dfm_1, sigmoid_table_784_4_sva_dfm_1,
          sigmoid_table_785_4_sva_dfm_1, sigmoid_table_786_4_sva_dfm_1, sigmoid_table_787_4_sva_dfm_1,
          sigmoid_table_788_4_sva_dfm_1, sigmoid_table_789_4_sva_dfm_1, sigmoid_table_790_4_sva_dfm_1,
          sigmoid_table_791_4_sva_dfm_1, sigmoid_table_792_4_sva_dfm_1, sigmoid_table_793_4_sva_dfm_1,
          sigmoid_table_794_4_sva_dfm_1, sigmoid_table_795_4_sva_dfm_1, sigmoid_table_796_4_sva_dfm_1,
          sigmoid_table_797_4_sva_dfm_1, sigmoid_table_798_4_sva_dfm_1, sigmoid_table_799_4_sva_dfm_1,
          sigmoid_table_800_4_sva_dfm_1, sigmoid_table_801_4_sva_dfm_1, sigmoid_table_802_4_sva_dfm_1,
          sigmoid_table_803_4_sva_dfm_1, sigmoid_table_804_4_sva_dfm_1, sigmoid_table_805_4_sva_dfm_1,
          sigmoid_table_806_4_sva_dfm_1, sigmoid_table_807_4_sva_dfm_1, sigmoid_table_808_4_sva_dfm_1,
          sigmoid_table_809_4_sva_dfm_1, sigmoid_table_810_4_sva_dfm_1, sigmoid_table_811_4_sva_dfm_1,
          sigmoid_table_812_4_sva_dfm_1, sigmoid_table_813_4_sva_dfm_1, sigmoid_table_814_4_sva_dfm_1,
          sigmoid_table_815_4_sva_dfm_1, sigmoid_table_816_4_sva_dfm_1, sigmoid_table_817_4_sva_dfm_1,
          sigmoid_table_818_4_sva_dfm_1, sigmoid_table_819_4_sva_dfm_1, sigmoid_table_820_4_sva_dfm_1,
          sigmoid_table_821_4_sva_dfm_1, sigmoid_table_822_3_sva_dfm_1, sigmoid_table_823_3_sva_dfm_1,
          sigmoid_table_824_3_sva_dfm_1, sigmoid_table_825_3_sva_dfm_1, sigmoid_table_826_3_sva_dfm_1,
          sigmoid_table_827_3_sva_dfm_1, sigmoid_table_828_3_sva_dfm_1, sigmoid_table_829_3_sva_dfm_1,
          sigmoid_table_830_3_sva_dfm_1, sigmoid_table_831_3_sva_dfm_1, sigmoid_table_832_3_sva_dfm_1,
          sigmoid_table_833_3_sva_dfm_1, sigmoid_table_834_3_sva_dfm_1, sigmoid_table_835_3_sva_dfm_1,
          sigmoid_table_836_3_sva_dfm_1, sigmoid_table_837_3_sva_dfm_1, sigmoid_table_838_3_sva_dfm_1,
          sigmoid_table_839_3_sva_dfm_1, sigmoid_table_840_3_sva_dfm_1, sigmoid_table_841_3_sva_dfm_1,
          sigmoid_table_842_3_sva_dfm_1, sigmoid_table_843_3_sva_dfm_1, sigmoid_table_844_3_sva_dfm_1,
          sigmoid_table_845_3_sva_dfm_1, sigmoid_table_846_3_sva_dfm_1, sigmoid_table_847_3_sva_dfm_1,
          sigmoid_table_848_3_sva_dfm_1, sigmoid_table_849_3_sva_dfm_1, sigmoid_table_850_3_sva_dfm_1,
          sigmoid_table_851_3_sva_dfm_1, sigmoid_table_852_3_sva_dfm_1, sigmoid_table_853_3_sva_dfm_1,
          sigmoid_table_854_3_sva_dfm_1, sigmoid_table_855_3_sva_dfm_1, sigmoid_table_856_3_sva_dfm_1,
          sigmoid_table_857_3_sva_dfm_1, sigmoid_table_858_3_sva_dfm_1, sigmoid_table_859_3_sva_dfm_1,
          sigmoid_table_860_3_sva_dfm_1, sigmoid_table_861_3_sva_dfm_1, sigmoid_table_862_3_sva_dfm_1,
          sigmoid_table_863_3_sva_dfm_1, sigmoid_table_864_3_sva_dfm_1, sigmoid_table_865_3_sva_dfm_1,
          sigmoid_table_866_3_sva_dfm_1, sigmoid_table_867_2_sva_dfm_1, sigmoid_table_868_2_sva_dfm_1,
          sigmoid_table_869_2_sva_dfm_1, sigmoid_table_870_2_sva_dfm_1, sigmoid_table_871_2_sva_dfm_1,
          sigmoid_table_872_2_sva_dfm_1, sigmoid_table_873_2_sva_dfm_1, sigmoid_table_874_2_sva_dfm_1,
          sigmoid_table_875_2_sva_dfm_1, sigmoid_table_876_2_sva_dfm_1, sigmoid_table_877_2_sva_dfm_1,
          sigmoid_table_878_2_sva_dfm_1, sigmoid_table_879_2_sva_dfm_1, sigmoid_table_880_2_sva_dfm_1,
          sigmoid_table_881_2_sva_dfm_1, sigmoid_table_882_2_sva_dfm_1, sigmoid_table_883_2_sva_dfm_1,
          sigmoid_table_884_2_sva_dfm_1, sigmoid_table_885_2_sva_dfm_1, sigmoid_table_886_2_sva_dfm_1,
          sigmoid_table_887_2_sva_dfm_1, sigmoid_table_888_2_sva_dfm_1, sigmoid_table_889_2_sva_dfm_1,
          sigmoid_table_890_2_sva_dfm_1, sigmoid_table_891_2_sva_dfm_1, sigmoid_table_892_2_sva_dfm_1,
          sigmoid_table_893_2_sva_dfm_1, sigmoid_table_894_2_sva_dfm_1, sigmoid_table_895_2_sva_dfm_1,
          sigmoid_table_896_2_sva_dfm_1, sigmoid_table_897_2_sva_dfm_1, sigmoid_table_898_2_sva_dfm_1,
          sigmoid_table_899_2_sva_dfm_1, sigmoid_table_900_2_sva_dfm_1, sigmoid_table_901_2_sva_dfm_1,
          sigmoid_table_902_2_sva_dfm_1, sigmoid_table_903_2_sva_dfm_1, sigmoid_table_904_2_sva_dfm_1,
          sigmoid_table_905_2_sva_dfm_1, sigmoid_table_906_2_sva_dfm_1, sigmoid_table_907_2_sva_dfm_1,
          sigmoid_table_908_2_sva_dfm_1, sigmoid_table_909_2_sva_dfm_1, sigmoid_table_910_2_sva_dfm_1,
          sigmoid_table_911_1_sva_dfm_1, sigmoid_table_912_1_sva_dfm_1, sigmoid_table_913_1_sva_dfm_1,
          sigmoid_table_914_1_sva_dfm_1, sigmoid_table_915_1_sva_dfm_1, sigmoid_table_916_1_sva_dfm_1,
          sigmoid_table_917_1_sva_dfm_1, sigmoid_table_918_1_sva_dfm_1, sigmoid_table_919_1_sva_dfm_1,
          sigmoid_table_920_1_sva_dfm_1, sigmoid_table_921_1_sva_dfm_1, sigmoid_table_922_1_sva_dfm_1,
          sigmoid_table_923_1_sva_dfm_1, sigmoid_table_924_1_sva_dfm_1, sigmoid_table_925_1_sva_dfm_1,
          sigmoid_table_926_1_sva_dfm_1, sigmoid_table_927_1_sva_dfm_1, sigmoid_table_928_1_sva_dfm_1,
          sigmoid_table_929_1_sva_dfm_1, sigmoid_table_930_1_sva_dfm_1, sigmoid_table_931_1_sva_dfm_1,
          sigmoid_table_932_1_sva_dfm_1, sigmoid_table_933_1_sva_dfm_1, sigmoid_table_934_1_sva_dfm_1,
          sigmoid_table_935_1_sva_dfm_1, sigmoid_table_936_1_sva_dfm_1, sigmoid_table_937_1_sva_dfm_1,
          sigmoid_table_938_1_sva_dfm_1, sigmoid_table_939_1_sva_dfm_1, sigmoid_table_940_1_sva_dfm_1,
          sigmoid_table_941_1_sva_dfm_1, sigmoid_table_942_1_sva_dfm_1, sigmoid_table_943_1_sva_dfm_1,
          sigmoid_table_944_1_sva_dfm_1, sigmoid_table_945_1_sva_dfm_1, sigmoid_table_946_1_sva_dfm_1,
          sigmoid_table_947_1_sva_dfm_1, sigmoid_table_948_1_sva_dfm_1, sigmoid_table_949_1_sva_dfm_1,
          sigmoid_table_950_1_sva_dfm_1, sigmoid_table_951_1_sva_dfm_1, sigmoid_table_952_1_sva_dfm_1,
          sigmoid_table_953_1_sva_dfm_1, sigmoid_table_954_1_sva_dfm_1, sigmoid_table_955_0_sva_dfm_1,
          sigmoid_table_956_0_sva_dfm_1, sigmoid_table_957_0_sva_dfm_1, sigmoid_table_958_0_sva_dfm_1,
          sigmoid_table_959_0_sva_dfm_1, sigmoid_table_960_0_sva_dfm_1, sigmoid_table_961_0_sva_dfm_1,
          sigmoid_table_962_0_sva_dfm_1, sigmoid_table_963_0_sva_dfm_1, sigmoid_table_964_0_sva_dfm_1,
          sigmoid_table_965_0_sva_dfm_1, sigmoid_table_966_0_sva_dfm_1, sigmoid_table_967_0_sva_dfm_1,
          sigmoid_table_968_0_sva_dfm_1, sigmoid_table_969_0_sva_dfm_1, sigmoid_table_970_0_sva_dfm_1,
          sigmoid_table_971_0_sva_dfm_1, sigmoid_table_972_0_sva_dfm_1, sigmoid_table_973_0_sva_dfm_1,
          sigmoid_table_974_0_sva_dfm_1, sigmoid_table_975_0_sva_dfm_1, sigmoid_table_976_0_sva_dfm_1,
          sigmoid_table_977_0_sva_dfm_1, sigmoid_table_978_0_sva_dfm_1, sigmoid_table_979_0_sva_dfm_1,
          sigmoid_table_980_0_sva_dfm_1, sigmoid_table_981_0_sva_dfm_1, sigmoid_table_982_0_sva_dfm_1,
          sigmoid_table_983_0_sva_dfm_1, sigmoid_table_984_0_sva_dfm_1, sigmoid_table_985_0_sva_dfm_1,
          sigmoid_table_986_0_sva_dfm_1, sigmoid_table_987_0_sva_dfm_1, sigmoid_table_988_0_sva_dfm_1,
          sigmoid_table_989_0_sva_dfm_1, sigmoid_table_990_0_sva_dfm_1, sigmoid_table_991_0_sva_dfm_1,
          sigmoid_table_992_0_sva_dfm_1, sigmoid_table_993_0_sva_dfm_1, sigmoid_table_994_0_sva_dfm_1,
          sigmoid_table_995_0_sva_dfm_1, sigmoid_table_996_0_sva_dfm_1, sigmoid_table_997_0_sva_dfm_1,
          sigmoid_table_998_0_sva_dfm_1, sigmoid_table_999_0_sva_dfm_1, sigmoid_table_1000_0_sva_dfm_1,
          sigmoid_table_1001_0_sva_dfm_1, sigmoid_table_1002_0_sva_dfm_1, sigmoid_table_1003_0_sva_dfm_1,
          sigmoid_table_1004_0_sva_dfm_1, sigmoid_table_1005_0_sva_dfm_1, sigmoid_table_1006_0_sva_dfm_1,
          sigmoid_table_1007_0_sva_dfm_1, sigmoid_table_1008_0_sva_dfm_1, sigmoid_table_1009_0_sva_dfm_1,
          sigmoid_table_1010_0_sva_dfm_1, sigmoid_table_1011_0_sva_dfm_1, sigmoid_table_1012_0_sva_dfm_1,
          sigmoid_table_1013_0_sva_dfm_1, sigmoid_table_1014_0_sva_dfm_1, sigmoid_table_1015_0_sva_dfm_1,
          sigmoid_table_1016_0_sva_dfm_1, sigmoid_table_1017_0_sva_dfm_1, sigmoid_table_1018_0_sva_dfm_1,
          sigmoid_table_1019_0_sva_dfm_1, sigmoid_table_1020_0_sva_dfm_1, sigmoid_table_1021_0_sva_dfm_1,
          sigmoid_table_1022_0_sva_dfm_1, sigmoid_table_1023_0_sva_dfm_1, {for_for_or_1_itm
          , for_for_or_itm});
      res_rsci_d_3 <= MUX_s_1_1024_2(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_202_3_sva_dfm_1, sigmoid_table_203_3_sva_dfm_1,
          sigmoid_table_204_3_sva_dfm_1, sigmoid_table_205_3_sva_dfm_1, sigmoid_table_206_3_sva_dfm_1,
          sigmoid_table_207_3_sva_dfm_1, sigmoid_table_208_3_sva_dfm_1, sigmoid_table_209_3_sva_dfm_1,
          sigmoid_table_210_3_sva_dfm_1, sigmoid_table_211_3_sva_dfm_1, sigmoid_table_212_3_sva_dfm_1,
          sigmoid_table_213_3_sva_dfm_1, sigmoid_table_214_3_sva_dfm_1, sigmoid_table_215_3_sva_dfm_1,
          sigmoid_table_216_3_sva_dfm_1, sigmoid_table_217_3_sva_dfm_1, sigmoid_table_218_3_sva_dfm_1,
          sigmoid_table_219_3_sva_dfm_1, sigmoid_table_220_3_sva_dfm_1, sigmoid_table_221_3_sva_dfm_1,
          sigmoid_table_222_3_sva_dfm_1, sigmoid_table_223_3_sva_dfm_1, sigmoid_table_224_3_sva_dfm_1,
          sigmoid_table_225_3_sva_dfm_1, sigmoid_table_226_3_sva_dfm_1, sigmoid_table_227_3_sva_dfm_1,
          sigmoid_table_228_3_sva_dfm_1, sigmoid_table_229_2_sva_dfm_1, sigmoid_table_230_2_sva_dfm_1,
          sigmoid_table_231_2_sva_dfm_1, sigmoid_table_232_2_sva_dfm_1, sigmoid_table_233_2_sva_dfm_1,
          sigmoid_table_234_2_sva_dfm_1, sigmoid_table_235_2_sva_dfm_1, sigmoid_table_236_2_sva_dfm_1,
          sigmoid_table_237_2_sva_dfm_1, sigmoid_table_238_2_sva_dfm_1, sigmoid_table_239_1_sva_dfm_1,
          sigmoid_table_240_1_sva_dfm_1, sigmoid_table_241_1_sva_dfm_1, sigmoid_table_242_1_sva_dfm_1,
          sigmoid_table_243_0_sva_dfm_1, sigmoid_table_244_0_sva_dfm_1, sigmoid_table_245_0_sva_dfm_1,
          sigmoid_table_246_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_274_3_sva_dfm_1,
          sigmoid_table_275_3_sva_dfm_1, sigmoid_table_276_3_sva_dfm_1, sigmoid_table_277_3_sva_dfm_1,
          sigmoid_table_278_3_sva_dfm_1, sigmoid_table_279_3_sva_dfm_1, sigmoid_table_280_3_sva_dfm_1,
          sigmoid_table_281_3_sva_dfm_1, sigmoid_table_282_3_sva_dfm_1, sigmoid_table_283_3_sva_dfm_1,
          sigmoid_table_284_2_sva_dfm_1, sigmoid_table_285_2_sva_dfm_1, sigmoid_table_286_2_sva_dfm_1,
          sigmoid_table_287_2_sva_dfm_1, sigmoid_table_288_1_sva_dfm_1, sigmoid_table_289_1_sva_dfm_1,
          sigmoid_table_290_1_sva_dfm_1, sigmoid_table_291_0_sva_dfm_1, sigmoid_table_292_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, sigmoid_table_308_3_sva_dfm_1, sigmoid_table_309_3_sva_dfm_1,
          sigmoid_table_310_3_sva_dfm_1, sigmoid_table_311_3_sva_dfm_1, sigmoid_table_312_3_sva_dfm_1,
          sigmoid_table_313_3_sva_dfm_1, sigmoid_table_314_2_sva_dfm_1, sigmoid_table_315_2_sva_dfm_1,
          sigmoid_table_316_2_sva_dfm_1, sigmoid_table_317_1_sva_dfm_1, sigmoid_table_318_0_sva_dfm_1,
          sigmoid_table_319_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, sigmoid_table_330_3_sva_dfm_1, sigmoid_table_331_3_sva_dfm_1,
          sigmoid_table_332_3_sva_dfm_1, sigmoid_table_333_3_sva_dfm_1, sigmoid_table_334_3_sva_dfm_1,
          sigmoid_table_335_2_sva_dfm_1, sigmoid_table_336_2_sva_dfm_1, sigmoid_table_337_1_sva_dfm_1,
          sigmoid_table_338_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, sigmoid_table_347_3_sva_dfm_1, sigmoid_table_348_3_sva_dfm_1, sigmoid_table_349_3_sva_dfm_1,
          sigmoid_table_350_3_sva_dfm_1, sigmoid_table_351_2_sva_dfm_1, sigmoid_table_352_2_sva_dfm_1,
          sigmoid_table_353_1_sva_dfm_1, sigmoid_table_354_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_361_3_sva_dfm_1, sigmoid_table_362_3_sva_dfm_1,
          sigmoid_table_363_3_sva_dfm_1, sigmoid_table_364_2_sva_dfm_1, sigmoid_table_365_2_sva_dfm_1,
          sigmoid_table_366_1_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_373_3_sva_dfm_1,
          sigmoid_table_374_3_sva_dfm_1, sigmoid_table_375_3_sva_dfm_1, sigmoid_table_376_2_sva_dfm_1,
          sigmoid_table_377_1_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_383_3_sva_dfm_1,
          sigmoid_table_384_3_sva_dfm_1, sigmoid_table_385_3_sva_dfm_1, sigmoid_table_386_2_sva_dfm_1,
          sigmoid_table_387_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_392_3_sva_dfm_1,
          sigmoid_table_393_3_sva_dfm_1, sigmoid_table_394_3_sva_dfm_1, sigmoid_table_395_2_sva_dfm_1,
          sigmoid_table_396_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_401_3_sva_dfm_1,
          sigmoid_table_402_3_sva_dfm_1, sigmoid_table_403_2_sva_dfm_1, sigmoid_table_404_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, sigmoid_table_408_3_sva_dfm_1, sigmoid_table_409_3_sva_dfm_1,
          sigmoid_table_410_2_sva_dfm_1, sigmoid_table_411_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, sigmoid_table_415_3_sva_dfm_1, sigmoid_table_416_3_sva_dfm_1, sigmoid_table_417_2_sva_dfm_1,
          sigmoid_table_418_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, sigmoid_table_422_3_sva_dfm_1,
          sigmoid_table_423_2_sva_dfm_1, sigmoid_table_424_1_sva_dfm_1, 1'b0, 1'b0,
          1'b0, sigmoid_table_428_3_sva_dfm_1, sigmoid_table_429_3_sva_dfm_1, sigmoid_table_430_1_sva_dfm_1,
          1'b0, 1'b0, 1'b0, sigmoid_table_434_3_sva_dfm_1, sigmoid_table_435_2_sva_dfm_1,
          sigmoid_table_436_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_439_3_sva_dfm_1,
          sigmoid_table_440_3_sva_dfm_1, sigmoid_table_441_2_sva_dfm_1, 1'b0, 1'b0,
          1'b0, sigmoid_table_445_3_sva_dfm_1, sigmoid_table_446_2_sva_dfm_1, 1'b0,
          1'b0, 1'b0, sigmoid_table_450_3_sva_dfm_1, sigmoid_table_451_2_sva_dfm_1,
          1'b0, 1'b0, 1'b0, sigmoid_table_455_3_sva_dfm_1, sigmoid_table_456_2_sva_dfm_1,
          1'b0, 1'b0, 1'b0, sigmoid_table_460_3_sva_dfm_1, sigmoid_table_461_1_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_464_3_sva_dfm_1, sigmoid_table_465_2_sva_dfm_1,
          sigmoid_table_466_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_469_3_sva_dfm_1,
          sigmoid_table_470_2_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_473_3_sva_dfm_1,
          sigmoid_table_474_2_sva_dfm_1, sigmoid_table_475_0_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_478_3_sva_dfm_1, sigmoid_table_479_1_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_482_3_sva_dfm_1, sigmoid_table_483_2_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_486_3_sva_dfm_1, sigmoid_table_487_2_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_490_3_sva_dfm_1, sigmoid_table_491_2_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_494_3_sva_dfm_1, sigmoid_table_495_2_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_498_3_sva_dfm_1, sigmoid_table_499_2_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_502_3_sva_dfm_1, sigmoid_table_503_2_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_506_3_sva_dfm_1, sigmoid_table_507_2_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_510_3_sva_dfm_1, sigmoid_table_511_2_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_514_3_sva_dfm_1, sigmoid_table_515_2_sva_dfm_1, sigmoid_table_516_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_519_3_sva_dfm_1, sigmoid_table_520_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_523_3_sva_dfm_1, sigmoid_table_524_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_527_3_sva_dfm_1, sigmoid_table_528_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_531_3_sva_dfm_1, sigmoid_table_532_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_535_3_sva_dfm_1, sigmoid_table_536_1_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_539_3_sva_dfm_1, sigmoid_table_540_1_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_543_3_sva_dfm_1, sigmoid_table_544_2_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_547_3_sva_dfm_1, sigmoid_table_548_2_sva_dfm_1,
          1'b0, 1'b0, 1'b0, sigmoid_table_552_3_sva_dfm_1, sigmoid_table_553_1_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_556_3_sva_dfm_1, sigmoid_table_557_2_sva_dfm_1,
          1'b0, 1'b0, 1'b0, sigmoid_table_561_3_sva_dfm_1, sigmoid_table_562_1_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_565_3_sva_dfm_1, sigmoid_table_566_2_sva_dfm_1,
          sigmoid_table_567_0_sva_dfm_1, 1'b0, 1'b0, sigmoid_table_570_3_sva_dfm_1,
          sigmoid_table_571_2_sva_dfm_1, sigmoid_table_572_0_sva_dfm_1, 1'b0, 1'b0,
          sigmoid_table_575_3_sva_dfm_1, sigmoid_table_576_2_sva_dfm_1, sigmoid_table_577_0_sva_dfm_1,
          1'b0, 1'b0, sigmoid_table_580_3_sva_dfm_1, sigmoid_table_581_2_sva_dfm_1,
          sigmoid_table_582_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, sigmoid_table_586_3_sva_dfm_1,
          sigmoid_table_587_2_sva_dfm_1, 1'b0, 1'b0, 1'b0, sigmoid_table_591_3_sva_dfm_1,
          sigmoid_table_592_3_sva_dfm_1, sigmoid_table_593_1_sva_dfm_1, 1'b0, 1'b0,
          1'b0, sigmoid_table_597_3_sva_dfm_1, sigmoid_table_598_2_sva_dfm_1, sigmoid_table_599_1_sva_dfm_1,
          1'b0, 1'b0, 1'b0, sigmoid_table_603_3_sva_dfm_1, sigmoid_table_604_3_sva_dfm_1,
          sigmoid_table_605_2_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_610_3_sva_dfm_1,
          sigmoid_table_611_2_sva_dfm_1, sigmoid_table_612_1_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_617_3_sva_dfm_1, sigmoid_table_618_3_sva_dfm_1,
          sigmoid_table_619_1_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_624_3_sva_dfm_1,
          sigmoid_table_625_3_sva_dfm_1, sigmoid_table_626_2_sva_dfm_1, sigmoid_table_627_1_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_633_3_sva_dfm_1, sigmoid_table_634_3_sva_dfm_1,
          sigmoid_table_635_2_sva_dfm_1, sigmoid_table_636_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, sigmoid_table_642_3_sva_dfm_1, sigmoid_table_643_3_sva_dfm_1,
          sigmoid_table_644_2_sva_dfm_1, sigmoid_table_645_1_sva_dfm_1, sigmoid_table_646_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_652_3_sva_dfm_1, sigmoid_table_653_3_sva_dfm_1,
          sigmoid_table_654_3_sva_dfm_1, sigmoid_table_655_2_sva_dfm_1, sigmoid_table_656_1_sva_dfm_1,
          sigmoid_table_657_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_664_3_sva_dfm_1,
          sigmoid_table_665_3_sva_dfm_1, sigmoid_table_666_3_sva_dfm_1, sigmoid_table_667_2_sva_dfm_1,
          sigmoid_table_668_2_sva_dfm_1, sigmoid_table_669_1_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_678_3_sva_dfm_1, sigmoid_table_679_3_sva_dfm_1,
          sigmoid_table_680_3_sva_dfm_1, sigmoid_table_681_3_sva_dfm_1, sigmoid_table_682_2_sva_dfm_1,
          sigmoid_table_683_2_sva_dfm_1, sigmoid_table_684_1_sva_dfm_1, sigmoid_table_685_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_695_3_sva_dfm_1,
          sigmoid_table_696_3_sva_dfm_1, sigmoid_table_697_3_sva_dfm_1, sigmoid_table_698_3_sva_dfm_1,
          sigmoid_table_699_3_sva_dfm_1, sigmoid_table_700_2_sva_dfm_1, sigmoid_table_701_2_sva_dfm_1,
          sigmoid_table_702_2_sva_dfm_1, sigmoid_table_703_1_sva_dfm_1, sigmoid_table_704_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          sigmoid_table_717_3_sva_dfm_1, sigmoid_table_718_3_sva_dfm_1, sigmoid_table_719_3_sva_dfm_1,
          sigmoid_table_720_3_sva_dfm_1, sigmoid_table_721_3_sva_dfm_1, sigmoid_table_722_3_sva_dfm_1,
          sigmoid_table_723_3_sva_dfm_1, sigmoid_table_724_2_sva_dfm_1, sigmoid_table_725_2_sva_dfm_1,
          sigmoid_table_726_2_sva_dfm_1, sigmoid_table_727_2_sva_dfm_1, sigmoid_table_728_1_sva_dfm_1,
          sigmoid_table_729_1_sva_dfm_1, sigmoid_table_730_0_sva_dfm_1, sigmoid_table_731_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_751_3_sva_dfm_1,
          sigmoid_table_752_3_sva_dfm_1, sigmoid_table_753_3_sva_dfm_1, sigmoid_table_754_3_sva_dfm_1,
          sigmoid_table_755_3_sva_dfm_1, sigmoid_table_756_3_sva_dfm_1, sigmoid_table_757_3_sva_dfm_1,
          sigmoid_table_758_3_sva_dfm_1, sigmoid_table_759_3_sva_dfm_1, sigmoid_table_760_3_sva_dfm_1,
          sigmoid_table_761_3_sva_dfm_1, sigmoid_table_762_3_sva_dfm_1, sigmoid_table_763_2_sva_dfm_1,
          sigmoid_table_764_2_sva_dfm_1, sigmoid_table_765_2_sva_dfm_1, sigmoid_table_766_2_sva_dfm_1,
          sigmoid_table_767_2_sva_dfm_1, sigmoid_table_768_2_sva_dfm_1, sigmoid_table_769_2_sva_dfm_1,
          sigmoid_table_770_1_sva_dfm_1, sigmoid_table_771_1_sva_dfm_1, sigmoid_table_772_1_sva_dfm_1,
          sigmoid_table_773_1_sva_dfm_1, sigmoid_table_774_0_sva_dfm_1, sigmoid_table_775_0_sva_dfm_1,
          sigmoid_table_776_0_sva_dfm_1, sigmoid_table_777_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_822_3_sva_dfm_1, sigmoid_table_823_3_sva_dfm_1,
          sigmoid_table_824_3_sva_dfm_1, sigmoid_table_825_3_sva_dfm_1, sigmoid_table_826_3_sva_dfm_1,
          sigmoid_table_827_3_sva_dfm_1, sigmoid_table_828_3_sva_dfm_1, sigmoid_table_829_3_sva_dfm_1,
          sigmoid_table_830_3_sva_dfm_1, sigmoid_table_831_3_sva_dfm_1, sigmoid_table_832_3_sva_dfm_1,
          sigmoid_table_833_3_sva_dfm_1, sigmoid_table_834_3_sva_dfm_1, sigmoid_table_835_3_sva_dfm_1,
          sigmoid_table_836_3_sva_dfm_1, sigmoid_table_837_3_sva_dfm_1, sigmoid_table_838_3_sva_dfm_1,
          sigmoid_table_839_3_sva_dfm_1, sigmoid_table_840_3_sva_dfm_1, sigmoid_table_841_3_sva_dfm_1,
          sigmoid_table_842_3_sva_dfm_1, sigmoid_table_843_3_sva_dfm_1, sigmoid_table_844_3_sva_dfm_1,
          sigmoid_table_845_3_sva_dfm_1, sigmoid_table_846_3_sva_dfm_1, sigmoid_table_847_3_sva_dfm_1,
          sigmoid_table_848_3_sva_dfm_1, sigmoid_table_849_3_sva_dfm_1, sigmoid_table_850_3_sva_dfm_1,
          sigmoid_table_851_3_sva_dfm_1, sigmoid_table_852_3_sva_dfm_1, sigmoid_table_853_3_sva_dfm_1,
          sigmoid_table_854_3_sva_dfm_1, sigmoid_table_855_3_sva_dfm_1, sigmoid_table_856_3_sva_dfm_1,
          sigmoid_table_857_3_sva_dfm_1, sigmoid_table_858_3_sva_dfm_1, sigmoid_table_859_3_sva_dfm_1,
          sigmoid_table_860_3_sva_dfm_1, sigmoid_table_861_3_sva_dfm_1, sigmoid_table_862_3_sva_dfm_1,
          sigmoid_table_863_3_sva_dfm_1, sigmoid_table_864_3_sva_dfm_1, sigmoid_table_865_3_sva_dfm_1,
          sigmoid_table_866_3_sva_dfm_1, sigmoid_table_867_2_sva_dfm_1, sigmoid_table_868_2_sva_dfm_1,
          sigmoid_table_869_2_sva_dfm_1, sigmoid_table_870_2_sva_dfm_1, sigmoid_table_871_2_sva_dfm_1,
          sigmoid_table_872_2_sva_dfm_1, sigmoid_table_873_2_sva_dfm_1, sigmoid_table_874_2_sva_dfm_1,
          sigmoid_table_875_2_sva_dfm_1, sigmoid_table_876_2_sva_dfm_1, sigmoid_table_877_2_sva_dfm_1,
          sigmoid_table_878_2_sva_dfm_1, sigmoid_table_879_2_sva_dfm_1, sigmoid_table_880_2_sva_dfm_1,
          sigmoid_table_881_2_sva_dfm_1, sigmoid_table_882_2_sva_dfm_1, sigmoid_table_883_2_sva_dfm_1,
          sigmoid_table_884_2_sva_dfm_1, sigmoid_table_885_2_sva_dfm_1, sigmoid_table_886_2_sva_dfm_1,
          sigmoid_table_887_2_sva_dfm_1, sigmoid_table_888_2_sva_dfm_1, sigmoid_table_889_2_sva_dfm_1,
          sigmoid_table_890_2_sva_dfm_1, sigmoid_table_891_2_sva_dfm_1, sigmoid_table_892_2_sva_dfm_1,
          sigmoid_table_893_2_sva_dfm_1, sigmoid_table_894_2_sva_dfm_1, sigmoid_table_895_2_sva_dfm_1,
          sigmoid_table_896_2_sva_dfm_1, sigmoid_table_897_2_sva_dfm_1, sigmoid_table_898_2_sva_dfm_1,
          sigmoid_table_899_2_sva_dfm_1, sigmoid_table_900_2_sva_dfm_1, sigmoid_table_901_2_sva_dfm_1,
          sigmoid_table_902_2_sva_dfm_1, sigmoid_table_903_2_sva_dfm_1, sigmoid_table_904_2_sva_dfm_1,
          sigmoid_table_905_2_sva_dfm_1, sigmoid_table_906_2_sva_dfm_1, sigmoid_table_907_2_sva_dfm_1,
          sigmoid_table_908_2_sva_dfm_1, sigmoid_table_909_2_sva_dfm_1, sigmoid_table_910_2_sva_dfm_1,
          sigmoid_table_911_1_sva_dfm_1, sigmoid_table_912_1_sva_dfm_1, sigmoid_table_913_1_sva_dfm_1,
          sigmoid_table_914_1_sva_dfm_1, sigmoid_table_915_1_sva_dfm_1, sigmoid_table_916_1_sva_dfm_1,
          sigmoid_table_917_1_sva_dfm_1, sigmoid_table_918_1_sva_dfm_1, sigmoid_table_919_1_sva_dfm_1,
          sigmoid_table_920_1_sva_dfm_1, sigmoid_table_921_1_sva_dfm_1, sigmoid_table_922_1_sva_dfm_1,
          sigmoid_table_923_1_sva_dfm_1, sigmoid_table_924_1_sva_dfm_1, sigmoid_table_925_1_sva_dfm_1,
          sigmoid_table_926_1_sva_dfm_1, sigmoid_table_927_1_sva_dfm_1, sigmoid_table_928_1_sva_dfm_1,
          sigmoid_table_929_1_sva_dfm_1, sigmoid_table_930_1_sva_dfm_1, sigmoid_table_931_1_sva_dfm_1,
          sigmoid_table_932_1_sva_dfm_1, sigmoid_table_933_1_sva_dfm_1, sigmoid_table_934_1_sva_dfm_1,
          sigmoid_table_935_1_sva_dfm_1, sigmoid_table_936_1_sva_dfm_1, sigmoid_table_937_1_sva_dfm_1,
          sigmoid_table_938_1_sva_dfm_1, sigmoid_table_939_1_sva_dfm_1, sigmoid_table_940_1_sva_dfm_1,
          sigmoid_table_941_1_sva_dfm_1, sigmoid_table_942_1_sva_dfm_1, sigmoid_table_943_1_sva_dfm_1,
          sigmoid_table_944_1_sva_dfm_1, sigmoid_table_945_1_sva_dfm_1, sigmoid_table_946_1_sva_dfm_1,
          sigmoid_table_947_1_sva_dfm_1, sigmoid_table_948_1_sva_dfm_1, sigmoid_table_949_1_sva_dfm_1,
          sigmoid_table_950_1_sva_dfm_1, sigmoid_table_951_1_sva_dfm_1, sigmoid_table_952_1_sva_dfm_1,
          sigmoid_table_953_1_sva_dfm_1, sigmoid_table_954_1_sva_dfm_1, sigmoid_table_955_0_sva_dfm_1,
          sigmoid_table_956_0_sva_dfm_1, sigmoid_table_957_0_sva_dfm_1, sigmoid_table_958_0_sva_dfm_1,
          sigmoid_table_959_0_sva_dfm_1, sigmoid_table_960_0_sva_dfm_1, sigmoid_table_961_0_sva_dfm_1,
          sigmoid_table_962_0_sva_dfm_1, sigmoid_table_963_0_sva_dfm_1, sigmoid_table_964_0_sva_dfm_1,
          sigmoid_table_965_0_sva_dfm_1, sigmoid_table_966_0_sva_dfm_1, sigmoid_table_967_0_sva_dfm_1,
          sigmoid_table_968_0_sva_dfm_1, sigmoid_table_969_0_sva_dfm_1, sigmoid_table_970_0_sva_dfm_1,
          sigmoid_table_971_0_sva_dfm_1, sigmoid_table_972_0_sva_dfm_1, sigmoid_table_973_0_sva_dfm_1,
          sigmoid_table_974_0_sva_dfm_1, sigmoid_table_975_0_sva_dfm_1, sigmoid_table_976_0_sva_dfm_1,
          sigmoid_table_977_0_sva_dfm_1, sigmoid_table_978_0_sva_dfm_1, sigmoid_table_979_0_sva_dfm_1,
          sigmoid_table_980_0_sva_dfm_1, sigmoid_table_981_0_sva_dfm_1, sigmoid_table_982_0_sva_dfm_1,
          sigmoid_table_983_0_sva_dfm_1, sigmoid_table_984_0_sva_dfm_1, sigmoid_table_985_0_sva_dfm_1,
          sigmoid_table_986_0_sva_dfm_1, sigmoid_table_987_0_sva_dfm_1, sigmoid_table_988_0_sva_dfm_1,
          sigmoid_table_989_0_sva_dfm_1, sigmoid_table_990_0_sva_dfm_1, sigmoid_table_991_0_sva_dfm_1,
          sigmoid_table_992_0_sva_dfm_1, sigmoid_table_993_0_sva_dfm_1, sigmoid_table_994_0_sva_dfm_1,
          sigmoid_table_995_0_sva_dfm_1, sigmoid_table_996_0_sva_dfm_1, sigmoid_table_997_0_sva_dfm_1,
          sigmoid_table_998_0_sva_dfm_1, sigmoid_table_999_0_sva_dfm_1, sigmoid_table_1000_0_sva_dfm_1,
          sigmoid_table_1001_0_sva_dfm_1, sigmoid_table_1002_0_sva_dfm_1, sigmoid_table_1003_0_sva_dfm_1,
          sigmoid_table_1004_0_sva_dfm_1, sigmoid_table_1005_0_sva_dfm_1, sigmoid_table_1006_0_sva_dfm_1,
          sigmoid_table_1007_0_sva_dfm_1, sigmoid_table_1008_0_sva_dfm_1, sigmoid_table_1009_0_sva_dfm_1,
          sigmoid_table_1010_0_sva_dfm_1, sigmoid_table_1011_0_sva_dfm_1, sigmoid_table_1012_0_sva_dfm_1,
          sigmoid_table_1013_0_sva_dfm_1, sigmoid_table_1014_0_sva_dfm_1, sigmoid_table_1015_0_sva_dfm_1,
          sigmoid_table_1016_0_sva_dfm_1, sigmoid_table_1017_0_sva_dfm_1, sigmoid_table_1018_0_sva_dfm_1,
          sigmoid_table_1019_0_sva_dfm_1, sigmoid_table_1020_0_sva_dfm_1, sigmoid_table_1021_0_sva_dfm_1,
          sigmoid_table_1022_0_sva_dfm_1, sigmoid_table_1023_0_sva_dfm_1, {for_for_or_1_itm
          , for_for_or_itm});
      res_rsci_d_6 <= MUX_s_1_1024_2(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_339_6_sva_dfm_1,
          sigmoid_table_340_6_sva_dfm_1, sigmoid_table_341_6_sva_dfm_1, sigmoid_table_342_6_sva_dfm_1,
          sigmoid_table_343_6_sva_dfm_1, sigmoid_table_344_6_sva_dfm_1, sigmoid_table_345_6_sva_dfm_1,
          sigmoid_table_346_6_sva_dfm_1, sigmoid_table_347_6_sva_dfm_1, sigmoid_table_348_6_sva_dfm_1,
          sigmoid_table_349_6_sva_dfm_1, sigmoid_table_350_6_sva_dfm_1, sigmoid_table_351_6_sva_dfm_1,
          sigmoid_table_352_6_sva_dfm_1, sigmoid_table_353_6_sva_dfm_1, sigmoid_table_354_6_sva_dfm_1,
          sigmoid_table_355_6_sva_dfm_1, sigmoid_table_356_6_sva_dfm_1, sigmoid_table_357_6_sva_dfm_1,
          sigmoid_table_358_6_sva_dfm_1, sigmoid_table_359_6_sva_dfm_1, sigmoid_table_360_6_sva_dfm_1,
          sigmoid_table_361_6_sva_dfm_1, sigmoid_table_362_6_sva_dfm_1, sigmoid_table_363_6_sva_dfm_1,
          sigmoid_table_364_6_sva_dfm_1, sigmoid_table_365_6_sva_dfm_1, sigmoid_table_366_6_sva_dfm_1,
          sigmoid_table_367_5_sva_dfm_1, sigmoid_table_368_5_sva_dfm_1, sigmoid_table_369_5_sva_dfm_1,
          sigmoid_table_370_5_sva_dfm_1, sigmoid_table_371_5_sva_dfm_1, sigmoid_table_372_5_sva_dfm_1,
          sigmoid_table_373_5_sva_dfm_1, sigmoid_table_374_5_sva_dfm_1, sigmoid_table_375_5_sva_dfm_1,
          sigmoid_table_376_5_sva_dfm_1, sigmoid_table_377_5_sva_dfm_1, sigmoid_table_378_4_sva_dfm_1,
          sigmoid_table_379_4_sva_dfm_1, sigmoid_table_380_4_sva_dfm_1, sigmoid_table_381_4_sva_dfm_1,
          sigmoid_table_382_4_sva_dfm_1, sigmoid_table_383_3_sva_dfm_1, sigmoid_table_384_3_sva_dfm_1,
          sigmoid_table_385_3_sva_dfm_1, sigmoid_table_386_2_sva_dfm_1, sigmoid_table_387_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_419_6_sva_dfm_1,
          sigmoid_table_420_6_sva_dfm_1, sigmoid_table_421_6_sva_dfm_1, sigmoid_table_422_6_sva_dfm_1,
          sigmoid_table_423_6_sva_dfm_1, sigmoid_table_424_6_sva_dfm_1, sigmoid_table_425_6_sva_dfm_1,
          sigmoid_table_426_6_sva_dfm_1, sigmoid_table_427_6_sva_dfm_1, sigmoid_table_428_6_sva_dfm_1,
          sigmoid_table_429_6_sva_dfm_1, sigmoid_table_430_6_sva_dfm_1, sigmoid_table_431_5_sva_dfm_1,
          sigmoid_table_432_5_sva_dfm_1, sigmoid_table_433_5_sva_dfm_1, sigmoid_table_434_5_sva_dfm_1,
          sigmoid_table_435_5_sva_dfm_1, sigmoid_table_436_5_sva_dfm_1, sigmoid_table_437_4_sva_dfm_1,
          sigmoid_table_438_4_sva_dfm_1, sigmoid_table_439_3_sva_dfm_1, sigmoid_table_440_3_sva_dfm_1,
          sigmoid_table_441_2_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, sigmoid_table_462_6_sva_dfm_1, sigmoid_table_463_6_sva_dfm_1, sigmoid_table_464_6_sva_dfm_1,
          sigmoid_table_465_6_sva_dfm_1, sigmoid_table_466_6_sva_dfm_1, sigmoid_table_467_6_sva_dfm_1,
          sigmoid_table_468_6_sva_dfm_1, sigmoid_table_469_6_sva_dfm_1, sigmoid_table_470_6_sva_dfm_1,
          sigmoid_table_471_5_sva_dfm_1, sigmoid_table_472_5_sva_dfm_1, sigmoid_table_473_5_sva_dfm_1,
          sigmoid_table_474_5_sva_dfm_1, sigmoid_table_475_5_sva_dfm_1, sigmoid_table_476_4_sva_dfm_1,
          sigmoid_table_477_4_sva_dfm_1, sigmoid_table_478_3_sva_dfm_1, sigmoid_table_479_1_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_496_6_sva_dfm_1, sigmoid_table_497_6_sva_dfm_1,
          sigmoid_table_498_6_sva_dfm_1, sigmoid_table_499_6_sva_dfm_1, sigmoid_table_500_6_sva_dfm_1,
          sigmoid_table_501_6_sva_dfm_1, sigmoid_table_502_6_sva_dfm_1, sigmoid_table_503_6_sva_dfm_1,
          sigmoid_table_504_5_sva_dfm_1, sigmoid_table_505_5_sva_dfm_1, sigmoid_table_506_5_sva_dfm_1,
          sigmoid_table_507_5_sva_dfm_1, sigmoid_table_508_4_sva_dfm_1, sigmoid_table_509_4_sva_dfm_1,
          sigmoid_table_510_3_sva_dfm_1, sigmoid_table_511_2_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, sigmoid_table_529_6_sva_dfm_1, sigmoid_table_530_6_sva_dfm_1,
          sigmoid_table_531_6_sva_dfm_1, sigmoid_table_532_6_sva_dfm_1, sigmoid_table_533_6_sva_dfm_1,
          sigmoid_table_534_6_sva_dfm_1, sigmoid_table_535_6_sva_dfm_1, sigmoid_table_536_6_sva_dfm_1,
          sigmoid_table_537_5_sva_dfm_1, sigmoid_table_538_5_sva_dfm_1, sigmoid_table_539_5_sva_dfm_1,
          sigmoid_table_540_5_sva_dfm_1, sigmoid_table_541_4_sva_dfm_1, sigmoid_table_542_4_sva_dfm_1,
          sigmoid_table_543_3_sva_dfm_1, sigmoid_table_544_2_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_563_6_sva_dfm_1, sigmoid_table_564_6_sva_dfm_1,
          sigmoid_table_565_6_sva_dfm_1, sigmoid_table_566_6_sva_dfm_1, sigmoid_table_567_6_sva_dfm_1,
          sigmoid_table_568_6_sva_dfm_1, sigmoid_table_569_6_sva_dfm_1, sigmoid_table_570_6_sva_dfm_1,
          sigmoid_table_571_6_sva_dfm_1, sigmoid_table_572_6_sva_dfm_1, sigmoid_table_573_5_sva_dfm_1,
          sigmoid_table_574_5_sva_dfm_1, sigmoid_table_575_5_sva_dfm_1, sigmoid_table_576_5_sva_dfm_1,
          sigmoid_table_577_5_sva_dfm_1, sigmoid_table_578_4_sva_dfm_1, sigmoid_table_579_4_sva_dfm_1,
          sigmoid_table_580_3_sva_dfm_1, sigmoid_table_581_2_sva_dfm_1, sigmoid_table_582_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_606_6_sva_dfm_1,
          sigmoid_table_607_6_sva_dfm_1, sigmoid_table_608_6_sva_dfm_1, sigmoid_table_609_6_sva_dfm_1,
          sigmoid_table_610_6_sva_dfm_1, sigmoid_table_611_6_sva_dfm_1, sigmoid_table_612_6_sva_dfm_1,
          sigmoid_table_613_6_sva_dfm_1, sigmoid_table_614_6_sva_dfm_1, sigmoid_table_615_6_sva_dfm_1,
          sigmoid_table_616_6_sva_dfm_1, sigmoid_table_617_6_sva_dfm_1, sigmoid_table_618_6_sva_dfm_1,
          sigmoid_table_619_6_sva_dfm_1, sigmoid_table_620_5_sva_dfm_1, sigmoid_table_621_5_sva_dfm_1,
          sigmoid_table_622_5_sva_dfm_1, sigmoid_table_623_5_sva_dfm_1, sigmoid_table_624_5_sva_dfm_1,
          sigmoid_table_625_5_sva_dfm_1, sigmoid_table_626_5_sva_dfm_1, sigmoid_table_627_5_sva_dfm_1,
          sigmoid_table_628_4_sva_dfm_1, sigmoid_table_629_4_sva_dfm_1, sigmoid_table_630_4_sva_dfm_1,
          sigmoid_table_631_4_sva_dfm_1, sigmoid_table_632_4_sva_dfm_1, sigmoid_table_633_3_sva_dfm_1,
          sigmoid_table_634_3_sva_dfm_1, sigmoid_table_635_2_sva_dfm_1, sigmoid_table_636_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, sigmoid_table_686_6_sva_dfm_1, sigmoid_table_687_6_sva_dfm_1, sigmoid_table_688_6_sva_dfm_1,
          sigmoid_table_689_6_sva_dfm_1, sigmoid_table_690_6_sva_dfm_1, sigmoid_table_691_6_sva_dfm_1,
          sigmoid_table_692_6_sva_dfm_1, sigmoid_table_693_6_sva_dfm_1, sigmoid_table_694_6_sva_dfm_1,
          sigmoid_table_695_6_sva_dfm_1, sigmoid_table_696_6_sva_dfm_1, sigmoid_table_697_6_sva_dfm_1,
          sigmoid_table_698_6_sva_dfm_1, sigmoid_table_699_6_sva_dfm_1, sigmoid_table_700_6_sva_dfm_1,
          sigmoid_table_701_6_sva_dfm_1, sigmoid_table_702_6_sva_dfm_1, sigmoid_table_703_6_sva_dfm_1,
          sigmoid_table_704_6_sva_dfm_1, sigmoid_table_705_6_sva_dfm_1, sigmoid_table_706_6_sva_dfm_1,
          sigmoid_table_707_6_sva_dfm_1, sigmoid_table_708_6_sva_dfm_1, sigmoid_table_709_6_sva_dfm_1,
          sigmoid_table_710_6_sva_dfm_1, sigmoid_table_711_6_sva_dfm_1, sigmoid_table_712_6_sva_dfm_1,
          sigmoid_table_713_6_sva_dfm_1, sigmoid_table_714_6_sva_dfm_1, sigmoid_table_715_6_sva_dfm_1,
          sigmoid_table_716_6_sva_dfm_1, sigmoid_table_717_6_sva_dfm_1, sigmoid_table_718_6_sva_dfm_1,
          sigmoid_table_719_6_sva_dfm_1, sigmoid_table_720_6_sva_dfm_1, sigmoid_table_721_6_sva_dfm_1,
          sigmoid_table_722_6_sva_dfm_1, sigmoid_table_723_6_sva_dfm_1, sigmoid_table_724_6_sva_dfm_1,
          sigmoid_table_725_6_sva_dfm_1, sigmoid_table_726_6_sva_dfm_1, sigmoid_table_727_6_sva_dfm_1,
          sigmoid_table_728_6_sva_dfm_1, sigmoid_table_729_6_sva_dfm_1, sigmoid_table_730_6_sva_dfm_1,
          sigmoid_table_731_6_sva_dfm_1, sigmoid_table_732_5_sva_dfm_1, sigmoid_table_733_5_sva_dfm_1,
          sigmoid_table_734_5_sva_dfm_1, sigmoid_table_735_5_sva_dfm_1, sigmoid_table_736_5_sva_dfm_1,
          sigmoid_table_737_5_sva_dfm_1, sigmoid_table_738_5_sva_dfm_1, sigmoid_table_739_5_sva_dfm_1,
          sigmoid_table_740_5_sva_dfm_1, sigmoid_table_741_5_sva_dfm_1, sigmoid_table_742_5_sva_dfm_1,
          sigmoid_table_743_5_sva_dfm_1, sigmoid_table_744_5_sva_dfm_1, sigmoid_table_745_5_sva_dfm_1,
          sigmoid_table_746_5_sva_dfm_1, sigmoid_table_747_5_sva_dfm_1, sigmoid_table_748_5_sva_dfm_1,
          sigmoid_table_749_5_sva_dfm_1, sigmoid_table_750_5_sva_dfm_1, sigmoid_table_751_5_sva_dfm_1,
          sigmoid_table_752_5_sva_dfm_1, sigmoid_table_753_5_sva_dfm_1, sigmoid_table_754_5_sva_dfm_1,
          sigmoid_table_755_5_sva_dfm_1, sigmoid_table_756_5_sva_dfm_1, sigmoid_table_757_5_sva_dfm_1,
          sigmoid_table_758_5_sva_dfm_1, sigmoid_table_759_5_sva_dfm_1, sigmoid_table_760_5_sva_dfm_1,
          sigmoid_table_761_5_sva_dfm_1, sigmoid_table_762_5_sva_dfm_1, sigmoid_table_763_5_sva_dfm_1,
          sigmoid_table_764_5_sva_dfm_1, sigmoid_table_765_5_sva_dfm_1, sigmoid_table_766_5_sva_dfm_1,
          sigmoid_table_767_5_sva_dfm_1, sigmoid_table_768_5_sva_dfm_1, sigmoid_table_769_5_sva_dfm_1,
          sigmoid_table_770_5_sva_dfm_1, sigmoid_table_771_5_sva_dfm_1, sigmoid_table_772_5_sva_dfm_1,
          sigmoid_table_773_5_sva_dfm_1, sigmoid_table_774_5_sva_dfm_1, sigmoid_table_775_5_sva_dfm_1,
          sigmoid_table_776_5_sva_dfm_1, sigmoid_table_777_5_sva_dfm_1, sigmoid_table_778_4_sva_dfm_1,
          sigmoid_table_779_4_sva_dfm_1, sigmoid_table_780_4_sva_dfm_1, sigmoid_table_781_4_sva_dfm_1,
          sigmoid_table_782_4_sva_dfm_1, sigmoid_table_783_4_sva_dfm_1, sigmoid_table_784_4_sva_dfm_1,
          sigmoid_table_785_4_sva_dfm_1, sigmoid_table_786_4_sva_dfm_1, sigmoid_table_787_4_sva_dfm_1,
          sigmoid_table_788_4_sva_dfm_1, sigmoid_table_789_4_sva_dfm_1, sigmoid_table_790_4_sva_dfm_1,
          sigmoid_table_791_4_sva_dfm_1, sigmoid_table_792_4_sva_dfm_1, sigmoid_table_793_4_sva_dfm_1,
          sigmoid_table_794_4_sva_dfm_1, sigmoid_table_795_4_sva_dfm_1, sigmoid_table_796_4_sva_dfm_1,
          sigmoid_table_797_4_sva_dfm_1, sigmoid_table_798_4_sva_dfm_1, sigmoid_table_799_4_sva_dfm_1,
          sigmoid_table_800_4_sva_dfm_1, sigmoid_table_801_4_sva_dfm_1, sigmoid_table_802_4_sva_dfm_1,
          sigmoid_table_803_4_sva_dfm_1, sigmoid_table_804_4_sva_dfm_1, sigmoid_table_805_4_sva_dfm_1,
          sigmoid_table_806_4_sva_dfm_1, sigmoid_table_807_4_sva_dfm_1, sigmoid_table_808_4_sva_dfm_1,
          sigmoid_table_809_4_sva_dfm_1, sigmoid_table_810_4_sva_dfm_1, sigmoid_table_811_4_sva_dfm_1,
          sigmoid_table_812_4_sva_dfm_1, sigmoid_table_813_4_sva_dfm_1, sigmoid_table_814_4_sva_dfm_1,
          sigmoid_table_815_4_sva_dfm_1, sigmoid_table_816_4_sva_dfm_1, sigmoid_table_817_4_sva_dfm_1,
          sigmoid_table_818_4_sva_dfm_1, sigmoid_table_819_4_sva_dfm_1, sigmoid_table_820_4_sva_dfm_1,
          sigmoid_table_821_4_sva_dfm_1, sigmoid_table_822_3_sva_dfm_1, sigmoid_table_823_3_sva_dfm_1,
          sigmoid_table_824_3_sva_dfm_1, sigmoid_table_825_3_sva_dfm_1, sigmoid_table_826_3_sva_dfm_1,
          sigmoid_table_827_3_sva_dfm_1, sigmoid_table_828_3_sva_dfm_1, sigmoid_table_829_3_sva_dfm_1,
          sigmoid_table_830_3_sva_dfm_1, sigmoid_table_831_3_sva_dfm_1, sigmoid_table_832_3_sva_dfm_1,
          sigmoid_table_833_3_sva_dfm_1, sigmoid_table_834_3_sva_dfm_1, sigmoid_table_835_3_sva_dfm_1,
          sigmoid_table_836_3_sva_dfm_1, sigmoid_table_837_3_sva_dfm_1, sigmoid_table_838_3_sva_dfm_1,
          sigmoid_table_839_3_sva_dfm_1, sigmoid_table_840_3_sva_dfm_1, sigmoid_table_841_3_sva_dfm_1,
          sigmoid_table_842_3_sva_dfm_1, sigmoid_table_843_3_sva_dfm_1, sigmoid_table_844_3_sva_dfm_1,
          sigmoid_table_845_3_sva_dfm_1, sigmoid_table_846_3_sva_dfm_1, sigmoid_table_847_3_sva_dfm_1,
          sigmoid_table_848_3_sva_dfm_1, sigmoid_table_849_3_sva_dfm_1, sigmoid_table_850_3_sva_dfm_1,
          sigmoid_table_851_3_sva_dfm_1, sigmoid_table_852_3_sva_dfm_1, sigmoid_table_853_3_sva_dfm_1,
          sigmoid_table_854_3_sva_dfm_1, sigmoid_table_855_3_sva_dfm_1, sigmoid_table_856_3_sva_dfm_1,
          sigmoid_table_857_3_sva_dfm_1, sigmoid_table_858_3_sva_dfm_1, sigmoid_table_859_3_sva_dfm_1,
          sigmoid_table_860_3_sva_dfm_1, sigmoid_table_861_3_sva_dfm_1, sigmoid_table_862_3_sva_dfm_1,
          sigmoid_table_863_3_sva_dfm_1, sigmoid_table_864_3_sva_dfm_1, sigmoid_table_865_3_sva_dfm_1,
          sigmoid_table_866_3_sva_dfm_1, sigmoid_table_867_2_sva_dfm_1, sigmoid_table_868_2_sva_dfm_1,
          sigmoid_table_869_2_sva_dfm_1, sigmoid_table_870_2_sva_dfm_1, sigmoid_table_871_2_sva_dfm_1,
          sigmoid_table_872_2_sva_dfm_1, sigmoid_table_873_2_sva_dfm_1, sigmoid_table_874_2_sva_dfm_1,
          sigmoid_table_875_2_sva_dfm_1, sigmoid_table_876_2_sva_dfm_1, sigmoid_table_877_2_sva_dfm_1,
          sigmoid_table_878_2_sva_dfm_1, sigmoid_table_879_2_sva_dfm_1, sigmoid_table_880_2_sva_dfm_1,
          sigmoid_table_881_2_sva_dfm_1, sigmoid_table_882_2_sva_dfm_1, sigmoid_table_883_2_sva_dfm_1,
          sigmoid_table_884_2_sva_dfm_1, sigmoid_table_885_2_sva_dfm_1, sigmoid_table_886_2_sva_dfm_1,
          sigmoid_table_887_2_sva_dfm_1, sigmoid_table_888_2_sva_dfm_1, sigmoid_table_889_2_sva_dfm_1,
          sigmoid_table_890_2_sva_dfm_1, sigmoid_table_891_2_sva_dfm_1, sigmoid_table_892_2_sva_dfm_1,
          sigmoid_table_893_2_sva_dfm_1, sigmoid_table_894_2_sva_dfm_1, sigmoid_table_895_2_sva_dfm_1,
          sigmoid_table_896_2_sva_dfm_1, sigmoid_table_897_2_sva_dfm_1, sigmoid_table_898_2_sva_dfm_1,
          sigmoid_table_899_2_sva_dfm_1, sigmoid_table_900_2_sva_dfm_1, sigmoid_table_901_2_sva_dfm_1,
          sigmoid_table_902_2_sva_dfm_1, sigmoid_table_903_2_sva_dfm_1, sigmoid_table_904_2_sva_dfm_1,
          sigmoid_table_905_2_sva_dfm_1, sigmoid_table_906_2_sva_dfm_1, sigmoid_table_907_2_sva_dfm_1,
          sigmoid_table_908_2_sva_dfm_1, sigmoid_table_909_2_sva_dfm_1, sigmoid_table_910_2_sva_dfm_1,
          sigmoid_table_911_1_sva_dfm_1, sigmoid_table_912_1_sva_dfm_1, sigmoid_table_913_1_sva_dfm_1,
          sigmoid_table_914_1_sva_dfm_1, sigmoid_table_915_1_sva_dfm_1, sigmoid_table_916_1_sva_dfm_1,
          sigmoid_table_917_1_sva_dfm_1, sigmoid_table_918_1_sva_dfm_1, sigmoid_table_919_1_sva_dfm_1,
          sigmoid_table_920_1_sva_dfm_1, sigmoid_table_921_1_sva_dfm_1, sigmoid_table_922_1_sva_dfm_1,
          sigmoid_table_923_1_sva_dfm_1, sigmoid_table_924_1_sva_dfm_1, sigmoid_table_925_1_sva_dfm_1,
          sigmoid_table_926_1_sva_dfm_1, sigmoid_table_927_1_sva_dfm_1, sigmoid_table_928_1_sva_dfm_1,
          sigmoid_table_929_1_sva_dfm_1, sigmoid_table_930_1_sva_dfm_1, sigmoid_table_931_1_sva_dfm_1,
          sigmoid_table_932_1_sva_dfm_1, sigmoid_table_933_1_sva_dfm_1, sigmoid_table_934_1_sva_dfm_1,
          sigmoid_table_935_1_sva_dfm_1, sigmoid_table_936_1_sva_dfm_1, sigmoid_table_937_1_sva_dfm_1,
          sigmoid_table_938_1_sva_dfm_1, sigmoid_table_939_1_sva_dfm_1, sigmoid_table_940_1_sva_dfm_1,
          sigmoid_table_941_1_sva_dfm_1, sigmoid_table_942_1_sva_dfm_1, sigmoid_table_943_1_sva_dfm_1,
          sigmoid_table_944_1_sva_dfm_1, sigmoid_table_945_1_sva_dfm_1, sigmoid_table_946_1_sva_dfm_1,
          sigmoid_table_947_1_sva_dfm_1, sigmoid_table_948_1_sva_dfm_1, sigmoid_table_949_1_sva_dfm_1,
          sigmoid_table_950_1_sva_dfm_1, sigmoid_table_951_1_sva_dfm_1, sigmoid_table_952_1_sva_dfm_1,
          sigmoid_table_953_1_sva_dfm_1, sigmoid_table_954_1_sva_dfm_1, sigmoid_table_955_0_sva_dfm_1,
          sigmoid_table_956_0_sva_dfm_1, sigmoid_table_957_0_sva_dfm_1, sigmoid_table_958_0_sva_dfm_1,
          sigmoid_table_959_0_sva_dfm_1, sigmoid_table_960_0_sva_dfm_1, sigmoid_table_961_0_sva_dfm_1,
          sigmoid_table_962_0_sva_dfm_1, sigmoid_table_963_0_sva_dfm_1, sigmoid_table_964_0_sva_dfm_1,
          sigmoid_table_965_0_sva_dfm_1, sigmoid_table_966_0_sva_dfm_1, sigmoid_table_967_0_sva_dfm_1,
          sigmoid_table_968_0_sva_dfm_1, sigmoid_table_969_0_sva_dfm_1, sigmoid_table_970_0_sva_dfm_1,
          sigmoid_table_971_0_sva_dfm_1, sigmoid_table_972_0_sva_dfm_1, sigmoid_table_973_0_sva_dfm_1,
          sigmoid_table_974_0_sva_dfm_1, sigmoid_table_975_0_sva_dfm_1, sigmoid_table_976_0_sva_dfm_1,
          sigmoid_table_977_0_sva_dfm_1, sigmoid_table_978_0_sva_dfm_1, sigmoid_table_979_0_sva_dfm_1,
          sigmoid_table_980_0_sva_dfm_1, sigmoid_table_981_0_sva_dfm_1, sigmoid_table_982_0_sva_dfm_1,
          sigmoid_table_983_0_sva_dfm_1, sigmoid_table_984_0_sva_dfm_1, sigmoid_table_985_0_sva_dfm_1,
          sigmoid_table_986_0_sva_dfm_1, sigmoid_table_987_0_sva_dfm_1, sigmoid_table_988_0_sva_dfm_1,
          sigmoid_table_989_0_sva_dfm_1, sigmoid_table_990_0_sva_dfm_1, sigmoid_table_991_0_sva_dfm_1,
          sigmoid_table_992_0_sva_dfm_1, sigmoid_table_993_0_sva_dfm_1, sigmoid_table_994_0_sva_dfm_1,
          sigmoid_table_995_0_sva_dfm_1, sigmoid_table_996_0_sva_dfm_1, sigmoid_table_997_0_sva_dfm_1,
          sigmoid_table_998_0_sva_dfm_1, sigmoid_table_999_0_sva_dfm_1, sigmoid_table_1000_0_sva_dfm_1,
          sigmoid_table_1001_0_sva_dfm_1, sigmoid_table_1002_0_sva_dfm_1, sigmoid_table_1003_0_sva_dfm_1,
          sigmoid_table_1004_0_sva_dfm_1, sigmoid_table_1005_0_sva_dfm_1, sigmoid_table_1006_0_sva_dfm_1,
          sigmoid_table_1007_0_sva_dfm_1, sigmoid_table_1008_0_sva_dfm_1, sigmoid_table_1009_0_sva_dfm_1,
          sigmoid_table_1010_0_sva_dfm_1, sigmoid_table_1011_0_sva_dfm_1, sigmoid_table_1012_0_sva_dfm_1,
          sigmoid_table_1013_0_sva_dfm_1, sigmoid_table_1014_0_sva_dfm_1, sigmoid_table_1015_0_sva_dfm_1,
          sigmoid_table_1016_0_sva_dfm_1, sigmoid_table_1017_0_sva_dfm_1, sigmoid_table_1018_0_sva_dfm_1,
          sigmoid_table_1019_0_sva_dfm_1, sigmoid_table_1020_0_sva_dfm_1, sigmoid_table_1021_0_sva_dfm_1,
          sigmoid_table_1022_0_sva_dfm_1, sigmoid_table_1023_0_sva_dfm_1, {for_for_or_1_itm
          , for_for_or_itm});
      res_rsci_d_4 <= MUX_s_1_1024_2(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_247_4_sva_dfm_1,
          sigmoid_table_248_4_sva_dfm_1, sigmoid_table_249_4_sva_dfm_1, sigmoid_table_250_4_sva_dfm_1,
          sigmoid_table_251_4_sva_dfm_1, sigmoid_table_252_4_sva_dfm_1, sigmoid_table_253_4_sva_dfm_1,
          sigmoid_table_254_4_sva_dfm_1, sigmoid_table_255_4_sva_dfm_1, sigmoid_table_256_4_sva_dfm_1,
          sigmoid_table_257_4_sva_dfm_1, sigmoid_table_258_4_sva_dfm_1, sigmoid_table_259_4_sva_dfm_1,
          sigmoid_table_260_4_sva_dfm_1, sigmoid_table_261_4_sva_dfm_1, sigmoid_table_262_4_sva_dfm_1,
          sigmoid_table_263_4_sva_dfm_1, sigmoid_table_264_4_sva_dfm_1, sigmoid_table_265_4_sva_dfm_1,
          sigmoid_table_266_4_sva_dfm_1, sigmoid_table_267_4_sva_dfm_1, sigmoid_table_268_4_sva_dfm_1,
          sigmoid_table_269_4_sva_dfm_1, sigmoid_table_270_4_sva_dfm_1, sigmoid_table_271_4_sva_dfm_1,
          sigmoid_table_272_4_sva_dfm_1, sigmoid_table_273_4_sva_dfm_1, sigmoid_table_274_3_sva_dfm_1,
          sigmoid_table_275_3_sva_dfm_1, sigmoid_table_276_3_sva_dfm_1, sigmoid_table_277_3_sva_dfm_1,
          sigmoid_table_278_3_sva_dfm_1, sigmoid_table_279_3_sva_dfm_1, sigmoid_table_280_3_sva_dfm_1,
          sigmoid_table_281_3_sva_dfm_1, sigmoid_table_282_3_sva_dfm_1, sigmoid_table_283_3_sva_dfm_1,
          sigmoid_table_284_2_sva_dfm_1, sigmoid_table_285_2_sva_dfm_1, sigmoid_table_286_2_sva_dfm_1,
          sigmoid_table_287_2_sva_dfm_1, sigmoid_table_288_1_sva_dfm_1, sigmoid_table_289_1_sva_dfm_1,
          sigmoid_table_290_1_sva_dfm_1, sigmoid_table_291_0_sva_dfm_1, sigmoid_table_292_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, sigmoid_table_320_4_sva_dfm_1, sigmoid_table_321_4_sva_dfm_1,
          sigmoid_table_322_4_sva_dfm_1, sigmoid_table_323_4_sva_dfm_1, sigmoid_table_324_4_sva_dfm_1,
          sigmoid_table_325_4_sva_dfm_1, sigmoid_table_326_4_sva_dfm_1, sigmoid_table_327_4_sva_dfm_1,
          sigmoid_table_328_4_sva_dfm_1, sigmoid_table_329_4_sva_dfm_1, sigmoid_table_330_3_sva_dfm_1,
          sigmoid_table_331_3_sva_dfm_1, sigmoid_table_332_3_sva_dfm_1, sigmoid_table_333_3_sva_dfm_1,
          sigmoid_table_334_3_sva_dfm_1, sigmoid_table_335_2_sva_dfm_1, sigmoid_table_336_2_sva_dfm_1,
          sigmoid_table_337_1_sva_dfm_1, sigmoid_table_338_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_355_4_sva_dfm_1, sigmoid_table_356_4_sva_dfm_1,
          sigmoid_table_357_4_sva_dfm_1, sigmoid_table_358_4_sva_dfm_1, sigmoid_table_359_4_sva_dfm_1,
          sigmoid_table_360_4_sva_dfm_1, sigmoid_table_361_3_sva_dfm_1, sigmoid_table_362_3_sva_dfm_1,
          sigmoid_table_363_3_sva_dfm_1, sigmoid_table_364_2_sva_dfm_1, sigmoid_table_365_2_sva_dfm_1,
          sigmoid_table_366_1_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_378_4_sva_dfm_1, sigmoid_table_379_4_sva_dfm_1,
          sigmoid_table_380_4_sva_dfm_1, sigmoid_table_381_4_sva_dfm_1, sigmoid_table_382_4_sva_dfm_1,
          sigmoid_table_383_3_sva_dfm_1, sigmoid_table_384_3_sva_dfm_1, sigmoid_table_385_3_sva_dfm_1,
          sigmoid_table_386_2_sva_dfm_1, sigmoid_table_387_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_397_4_sva_dfm_1,
          sigmoid_table_398_4_sva_dfm_1, sigmoid_table_399_4_sva_dfm_1, sigmoid_table_400_4_sva_dfm_1,
          sigmoid_table_401_3_sva_dfm_1, sigmoid_table_402_3_sva_dfm_1, sigmoid_table_403_2_sva_dfm_1,
          sigmoid_table_404_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          sigmoid_table_412_4_sva_dfm_1, sigmoid_table_413_4_sva_dfm_1, sigmoid_table_414_4_sva_dfm_1,
          sigmoid_table_415_3_sva_dfm_1, sigmoid_table_416_3_sva_dfm_1, sigmoid_table_417_2_sva_dfm_1,
          sigmoid_table_418_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_425_4_sva_dfm_1,
          sigmoid_table_426_4_sva_dfm_1, sigmoid_table_427_4_sva_dfm_1, sigmoid_table_428_3_sva_dfm_1,
          sigmoid_table_429_3_sva_dfm_1, sigmoid_table_430_1_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_437_4_sva_dfm_1, sigmoid_table_438_4_sva_dfm_1,
          sigmoid_table_439_3_sva_dfm_1, sigmoid_table_440_3_sva_dfm_1, sigmoid_table_441_2_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_447_4_sva_dfm_1, sigmoid_table_448_4_sva_dfm_1,
          sigmoid_table_449_4_sva_dfm_1, sigmoid_table_450_3_sva_dfm_1, sigmoid_table_451_2_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_457_4_sva_dfm_1, sigmoid_table_458_4_sva_dfm_1,
          sigmoid_table_459_4_sva_dfm_1, sigmoid_table_460_3_sva_dfm_1, sigmoid_table_461_1_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_467_4_sva_dfm_1, sigmoid_table_468_4_sva_dfm_1,
          sigmoid_table_469_3_sva_dfm_1, sigmoid_table_470_2_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, sigmoid_table_476_4_sva_dfm_1, sigmoid_table_477_4_sva_dfm_1,
          sigmoid_table_478_3_sva_dfm_1, sigmoid_table_479_1_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_484_4_sva_dfm_1, sigmoid_table_485_4_sva_dfm_1,
          sigmoid_table_486_3_sva_dfm_1, sigmoid_table_487_2_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_492_4_sva_dfm_1, sigmoid_table_493_4_sva_dfm_1,
          sigmoid_table_494_3_sva_dfm_1, sigmoid_table_495_2_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_500_4_sva_dfm_1, sigmoid_table_501_4_sva_dfm_1,
          sigmoid_table_502_3_sva_dfm_1, sigmoid_table_503_2_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_508_4_sva_dfm_1, sigmoid_table_509_4_sva_dfm_1,
          sigmoid_table_510_3_sva_dfm_1, sigmoid_table_511_2_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, sigmoid_table_517_4_sva_dfm_1, sigmoid_table_518_4_sva_dfm_1,
          sigmoid_table_519_3_sva_dfm_1, sigmoid_table_520_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_525_4_sva_dfm_1, sigmoid_table_526_4_sva_dfm_1,
          sigmoid_table_527_3_sva_dfm_1, sigmoid_table_528_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_533_4_sva_dfm_1, sigmoid_table_534_4_sva_dfm_1,
          sigmoid_table_535_3_sva_dfm_1, sigmoid_table_536_1_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_541_4_sva_dfm_1, sigmoid_table_542_4_sva_dfm_1,
          sigmoid_table_543_3_sva_dfm_1, sigmoid_table_544_2_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_549_4_sva_dfm_1, sigmoid_table_550_4_sva_dfm_1,
          sigmoid_table_551_4_sva_dfm_1, sigmoid_table_552_3_sva_dfm_1, sigmoid_table_553_1_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_558_4_sva_dfm_1, sigmoid_table_559_4_sva_dfm_1,
          sigmoid_table_560_4_sva_dfm_1, sigmoid_table_561_3_sva_dfm_1, sigmoid_table_562_1_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_568_4_sva_dfm_1, sigmoid_table_569_4_sva_dfm_1,
          sigmoid_table_570_3_sva_dfm_1, sigmoid_table_571_2_sva_dfm_1, sigmoid_table_572_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_578_4_sva_dfm_1, sigmoid_table_579_4_sva_dfm_1,
          sigmoid_table_580_3_sva_dfm_1, sigmoid_table_581_2_sva_dfm_1, sigmoid_table_582_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_588_4_sva_dfm_1, sigmoid_table_589_4_sva_dfm_1,
          sigmoid_table_590_4_sva_dfm_1, sigmoid_table_591_3_sva_dfm_1, sigmoid_table_592_3_sva_dfm_1,
          sigmoid_table_593_1_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_600_4_sva_dfm_1,
          sigmoid_table_601_4_sva_dfm_1, sigmoid_table_602_4_sva_dfm_1, sigmoid_table_603_3_sva_dfm_1,
          sigmoid_table_604_3_sva_dfm_1, sigmoid_table_605_2_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_613_4_sva_dfm_1, sigmoid_table_614_4_sva_dfm_1,
          sigmoid_table_615_4_sva_dfm_1, sigmoid_table_616_4_sva_dfm_1, sigmoid_table_617_3_sva_dfm_1,
          sigmoid_table_618_3_sva_dfm_1, sigmoid_table_619_1_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_628_4_sva_dfm_1, sigmoid_table_629_4_sva_dfm_1,
          sigmoid_table_630_4_sva_dfm_1, sigmoid_table_631_4_sva_dfm_1, sigmoid_table_632_4_sva_dfm_1,
          sigmoid_table_633_3_sva_dfm_1, sigmoid_table_634_3_sva_dfm_1, sigmoid_table_635_2_sva_dfm_1,
          sigmoid_table_636_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, sigmoid_table_647_4_sva_dfm_1, sigmoid_table_648_4_sva_dfm_1,
          sigmoid_table_649_4_sva_dfm_1, sigmoid_table_650_4_sva_dfm_1, sigmoid_table_651_4_sva_dfm_1,
          sigmoid_table_652_3_sva_dfm_1, sigmoid_table_653_3_sva_dfm_1, sigmoid_table_654_3_sva_dfm_1,
          sigmoid_table_655_2_sva_dfm_1, sigmoid_table_656_1_sva_dfm_1, sigmoid_table_657_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          sigmoid_table_670_4_sva_dfm_1, sigmoid_table_671_4_sva_dfm_1, sigmoid_table_672_4_sva_dfm_1,
          sigmoid_table_673_4_sva_dfm_1, sigmoid_table_674_4_sva_dfm_1, sigmoid_table_675_4_sva_dfm_1,
          sigmoid_table_676_4_sva_dfm_1, sigmoid_table_677_4_sva_dfm_1, sigmoid_table_678_3_sva_dfm_1,
          sigmoid_table_679_3_sva_dfm_1, sigmoid_table_680_3_sva_dfm_1, sigmoid_table_681_3_sva_dfm_1,
          sigmoid_table_682_2_sva_dfm_1, sigmoid_table_683_2_sva_dfm_1, sigmoid_table_684_1_sva_dfm_1,
          sigmoid_table_685_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          sigmoid_table_705_4_sva_dfm_1, sigmoid_table_706_4_sva_dfm_1, sigmoid_table_707_4_sva_dfm_1,
          sigmoid_table_708_4_sva_dfm_1, sigmoid_table_709_4_sva_dfm_1, sigmoid_table_710_4_sva_dfm_1,
          sigmoid_table_711_4_sva_dfm_1, sigmoid_table_712_4_sva_dfm_1, sigmoid_table_713_4_sva_dfm_1,
          sigmoid_table_714_4_sva_dfm_1, sigmoid_table_715_4_sva_dfm_1, sigmoid_table_716_4_sva_dfm_1,
          sigmoid_table_717_3_sva_dfm_1, sigmoid_table_718_3_sva_dfm_1, sigmoid_table_719_3_sva_dfm_1,
          sigmoid_table_720_3_sva_dfm_1, sigmoid_table_721_3_sva_dfm_1, sigmoid_table_722_3_sva_dfm_1,
          sigmoid_table_723_3_sva_dfm_1, sigmoid_table_724_2_sva_dfm_1, sigmoid_table_725_2_sva_dfm_1,
          sigmoid_table_726_2_sva_dfm_1, sigmoid_table_727_2_sva_dfm_1, sigmoid_table_728_1_sva_dfm_1,
          sigmoid_table_729_1_sva_dfm_1, sigmoid_table_730_0_sva_dfm_1, sigmoid_table_731_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_778_4_sva_dfm_1,
          sigmoid_table_779_4_sva_dfm_1, sigmoid_table_780_4_sva_dfm_1, sigmoid_table_781_4_sva_dfm_1,
          sigmoid_table_782_4_sva_dfm_1, sigmoid_table_783_4_sva_dfm_1, sigmoid_table_784_4_sva_dfm_1,
          sigmoid_table_785_4_sva_dfm_1, sigmoid_table_786_4_sva_dfm_1, sigmoid_table_787_4_sva_dfm_1,
          sigmoid_table_788_4_sva_dfm_1, sigmoid_table_789_4_sva_dfm_1, sigmoid_table_790_4_sva_dfm_1,
          sigmoid_table_791_4_sva_dfm_1, sigmoid_table_792_4_sva_dfm_1, sigmoid_table_793_4_sva_dfm_1,
          sigmoid_table_794_4_sva_dfm_1, sigmoid_table_795_4_sva_dfm_1, sigmoid_table_796_4_sva_dfm_1,
          sigmoid_table_797_4_sva_dfm_1, sigmoid_table_798_4_sva_dfm_1, sigmoid_table_799_4_sva_dfm_1,
          sigmoid_table_800_4_sva_dfm_1, sigmoid_table_801_4_sva_dfm_1, sigmoid_table_802_4_sva_dfm_1,
          sigmoid_table_803_4_sva_dfm_1, sigmoid_table_804_4_sva_dfm_1, sigmoid_table_805_4_sva_dfm_1,
          sigmoid_table_806_4_sva_dfm_1, sigmoid_table_807_4_sva_dfm_1, sigmoid_table_808_4_sva_dfm_1,
          sigmoid_table_809_4_sva_dfm_1, sigmoid_table_810_4_sva_dfm_1, sigmoid_table_811_4_sva_dfm_1,
          sigmoid_table_812_4_sva_dfm_1, sigmoid_table_813_4_sva_dfm_1, sigmoid_table_814_4_sva_dfm_1,
          sigmoid_table_815_4_sva_dfm_1, sigmoid_table_816_4_sva_dfm_1, sigmoid_table_817_4_sva_dfm_1,
          sigmoid_table_818_4_sva_dfm_1, sigmoid_table_819_4_sva_dfm_1, sigmoid_table_820_4_sva_dfm_1,
          sigmoid_table_821_4_sva_dfm_1, sigmoid_table_822_3_sva_dfm_1, sigmoid_table_823_3_sva_dfm_1,
          sigmoid_table_824_3_sva_dfm_1, sigmoid_table_825_3_sva_dfm_1, sigmoid_table_826_3_sva_dfm_1,
          sigmoid_table_827_3_sva_dfm_1, sigmoid_table_828_3_sva_dfm_1, sigmoid_table_829_3_sva_dfm_1,
          sigmoid_table_830_3_sva_dfm_1, sigmoid_table_831_3_sva_dfm_1, sigmoid_table_832_3_sva_dfm_1,
          sigmoid_table_833_3_sva_dfm_1, sigmoid_table_834_3_sva_dfm_1, sigmoid_table_835_3_sva_dfm_1,
          sigmoid_table_836_3_sva_dfm_1, sigmoid_table_837_3_sva_dfm_1, sigmoid_table_838_3_sva_dfm_1,
          sigmoid_table_839_3_sva_dfm_1, sigmoid_table_840_3_sva_dfm_1, sigmoid_table_841_3_sva_dfm_1,
          sigmoid_table_842_3_sva_dfm_1, sigmoid_table_843_3_sva_dfm_1, sigmoid_table_844_3_sva_dfm_1,
          sigmoid_table_845_3_sva_dfm_1, sigmoid_table_846_3_sva_dfm_1, sigmoid_table_847_3_sva_dfm_1,
          sigmoid_table_848_3_sva_dfm_1, sigmoid_table_849_3_sva_dfm_1, sigmoid_table_850_3_sva_dfm_1,
          sigmoid_table_851_3_sva_dfm_1, sigmoid_table_852_3_sva_dfm_1, sigmoid_table_853_3_sva_dfm_1,
          sigmoid_table_854_3_sva_dfm_1, sigmoid_table_855_3_sva_dfm_1, sigmoid_table_856_3_sva_dfm_1,
          sigmoid_table_857_3_sva_dfm_1, sigmoid_table_858_3_sva_dfm_1, sigmoid_table_859_3_sva_dfm_1,
          sigmoid_table_860_3_sva_dfm_1, sigmoid_table_861_3_sva_dfm_1, sigmoid_table_862_3_sva_dfm_1,
          sigmoid_table_863_3_sva_dfm_1, sigmoid_table_864_3_sva_dfm_1, sigmoid_table_865_3_sva_dfm_1,
          sigmoid_table_866_3_sva_dfm_1, sigmoid_table_867_2_sva_dfm_1, sigmoid_table_868_2_sva_dfm_1,
          sigmoid_table_869_2_sva_dfm_1, sigmoid_table_870_2_sva_dfm_1, sigmoid_table_871_2_sva_dfm_1,
          sigmoid_table_872_2_sva_dfm_1, sigmoid_table_873_2_sva_dfm_1, sigmoid_table_874_2_sva_dfm_1,
          sigmoid_table_875_2_sva_dfm_1, sigmoid_table_876_2_sva_dfm_1, sigmoid_table_877_2_sva_dfm_1,
          sigmoid_table_878_2_sva_dfm_1, sigmoid_table_879_2_sva_dfm_1, sigmoid_table_880_2_sva_dfm_1,
          sigmoid_table_881_2_sva_dfm_1, sigmoid_table_882_2_sva_dfm_1, sigmoid_table_883_2_sva_dfm_1,
          sigmoid_table_884_2_sva_dfm_1, sigmoid_table_885_2_sva_dfm_1, sigmoid_table_886_2_sva_dfm_1,
          sigmoid_table_887_2_sva_dfm_1, sigmoid_table_888_2_sva_dfm_1, sigmoid_table_889_2_sva_dfm_1,
          sigmoid_table_890_2_sva_dfm_1, sigmoid_table_891_2_sva_dfm_1, sigmoid_table_892_2_sva_dfm_1,
          sigmoid_table_893_2_sva_dfm_1, sigmoid_table_894_2_sva_dfm_1, sigmoid_table_895_2_sva_dfm_1,
          sigmoid_table_896_2_sva_dfm_1, sigmoid_table_897_2_sva_dfm_1, sigmoid_table_898_2_sva_dfm_1,
          sigmoid_table_899_2_sva_dfm_1, sigmoid_table_900_2_sva_dfm_1, sigmoid_table_901_2_sva_dfm_1,
          sigmoid_table_902_2_sva_dfm_1, sigmoid_table_903_2_sva_dfm_1, sigmoid_table_904_2_sva_dfm_1,
          sigmoid_table_905_2_sva_dfm_1, sigmoid_table_906_2_sva_dfm_1, sigmoid_table_907_2_sva_dfm_1,
          sigmoid_table_908_2_sva_dfm_1, sigmoid_table_909_2_sva_dfm_1, sigmoid_table_910_2_sva_dfm_1,
          sigmoid_table_911_1_sva_dfm_1, sigmoid_table_912_1_sva_dfm_1, sigmoid_table_913_1_sva_dfm_1,
          sigmoid_table_914_1_sva_dfm_1, sigmoid_table_915_1_sva_dfm_1, sigmoid_table_916_1_sva_dfm_1,
          sigmoid_table_917_1_sva_dfm_1, sigmoid_table_918_1_sva_dfm_1, sigmoid_table_919_1_sva_dfm_1,
          sigmoid_table_920_1_sva_dfm_1, sigmoid_table_921_1_sva_dfm_1, sigmoid_table_922_1_sva_dfm_1,
          sigmoid_table_923_1_sva_dfm_1, sigmoid_table_924_1_sva_dfm_1, sigmoid_table_925_1_sva_dfm_1,
          sigmoid_table_926_1_sva_dfm_1, sigmoid_table_927_1_sva_dfm_1, sigmoid_table_928_1_sva_dfm_1,
          sigmoid_table_929_1_sva_dfm_1, sigmoid_table_930_1_sva_dfm_1, sigmoid_table_931_1_sva_dfm_1,
          sigmoid_table_932_1_sva_dfm_1, sigmoid_table_933_1_sva_dfm_1, sigmoid_table_934_1_sva_dfm_1,
          sigmoid_table_935_1_sva_dfm_1, sigmoid_table_936_1_sva_dfm_1, sigmoid_table_937_1_sva_dfm_1,
          sigmoid_table_938_1_sva_dfm_1, sigmoid_table_939_1_sva_dfm_1, sigmoid_table_940_1_sva_dfm_1,
          sigmoid_table_941_1_sva_dfm_1, sigmoid_table_942_1_sva_dfm_1, sigmoid_table_943_1_sva_dfm_1,
          sigmoid_table_944_1_sva_dfm_1, sigmoid_table_945_1_sva_dfm_1, sigmoid_table_946_1_sva_dfm_1,
          sigmoid_table_947_1_sva_dfm_1, sigmoid_table_948_1_sva_dfm_1, sigmoid_table_949_1_sva_dfm_1,
          sigmoid_table_950_1_sva_dfm_1, sigmoid_table_951_1_sva_dfm_1, sigmoid_table_952_1_sva_dfm_1,
          sigmoid_table_953_1_sva_dfm_1, sigmoid_table_954_1_sva_dfm_1, sigmoid_table_955_0_sva_dfm_1,
          sigmoid_table_956_0_sva_dfm_1, sigmoid_table_957_0_sva_dfm_1, sigmoid_table_958_0_sva_dfm_1,
          sigmoid_table_959_0_sva_dfm_1, sigmoid_table_960_0_sva_dfm_1, sigmoid_table_961_0_sva_dfm_1,
          sigmoid_table_962_0_sva_dfm_1, sigmoid_table_963_0_sva_dfm_1, sigmoid_table_964_0_sva_dfm_1,
          sigmoid_table_965_0_sva_dfm_1, sigmoid_table_966_0_sva_dfm_1, sigmoid_table_967_0_sva_dfm_1,
          sigmoid_table_968_0_sva_dfm_1, sigmoid_table_969_0_sva_dfm_1, sigmoid_table_970_0_sva_dfm_1,
          sigmoid_table_971_0_sva_dfm_1, sigmoid_table_972_0_sva_dfm_1, sigmoid_table_973_0_sva_dfm_1,
          sigmoid_table_974_0_sva_dfm_1, sigmoid_table_975_0_sva_dfm_1, sigmoid_table_976_0_sva_dfm_1,
          sigmoid_table_977_0_sva_dfm_1, sigmoid_table_978_0_sva_dfm_1, sigmoid_table_979_0_sva_dfm_1,
          sigmoid_table_980_0_sva_dfm_1, sigmoid_table_981_0_sva_dfm_1, sigmoid_table_982_0_sva_dfm_1,
          sigmoid_table_983_0_sva_dfm_1, sigmoid_table_984_0_sva_dfm_1, sigmoid_table_985_0_sva_dfm_1,
          sigmoid_table_986_0_sva_dfm_1, sigmoid_table_987_0_sva_dfm_1, sigmoid_table_988_0_sva_dfm_1,
          sigmoid_table_989_0_sva_dfm_1, sigmoid_table_990_0_sva_dfm_1, sigmoid_table_991_0_sva_dfm_1,
          sigmoid_table_992_0_sva_dfm_1, sigmoid_table_993_0_sva_dfm_1, sigmoid_table_994_0_sva_dfm_1,
          sigmoid_table_995_0_sva_dfm_1, sigmoid_table_996_0_sva_dfm_1, sigmoid_table_997_0_sva_dfm_1,
          sigmoid_table_998_0_sva_dfm_1, sigmoid_table_999_0_sva_dfm_1, sigmoid_table_1000_0_sva_dfm_1,
          sigmoid_table_1001_0_sva_dfm_1, sigmoid_table_1002_0_sva_dfm_1, sigmoid_table_1003_0_sva_dfm_1,
          sigmoid_table_1004_0_sva_dfm_1, sigmoid_table_1005_0_sva_dfm_1, sigmoid_table_1006_0_sva_dfm_1,
          sigmoid_table_1007_0_sva_dfm_1, sigmoid_table_1008_0_sva_dfm_1, sigmoid_table_1009_0_sva_dfm_1,
          sigmoid_table_1010_0_sva_dfm_1, sigmoid_table_1011_0_sva_dfm_1, sigmoid_table_1012_0_sva_dfm_1,
          sigmoid_table_1013_0_sva_dfm_1, sigmoid_table_1014_0_sva_dfm_1, sigmoid_table_1015_0_sva_dfm_1,
          sigmoid_table_1016_0_sva_dfm_1, sigmoid_table_1017_0_sva_dfm_1, sigmoid_table_1018_0_sva_dfm_1,
          sigmoid_table_1019_0_sva_dfm_1, sigmoid_table_1020_0_sva_dfm_1, sigmoid_table_1021_0_sva_dfm_1,
          sigmoid_table_1022_0_sva_dfm_1, sigmoid_table_1023_0_sva_dfm_1, {for_for_or_1_itm
          , for_for_or_itm});
      res_rsci_d_5 <= MUX_s_1_1024_2(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_293_5_sva_dfm_1,
          sigmoid_table_294_5_sva_dfm_1, sigmoid_table_295_5_sva_dfm_1, sigmoid_table_296_5_sva_dfm_1,
          sigmoid_table_297_5_sva_dfm_1, sigmoid_table_298_5_sva_dfm_1, sigmoid_table_299_5_sva_dfm_1,
          sigmoid_table_300_5_sva_dfm_1, sigmoid_table_301_5_sva_dfm_1, sigmoid_table_302_5_sva_dfm_1,
          sigmoid_table_303_5_sva_dfm_1, sigmoid_table_304_5_sva_dfm_1, sigmoid_table_305_5_sva_dfm_1,
          sigmoid_table_306_5_sva_dfm_1, sigmoid_table_307_5_sva_dfm_1, sigmoid_table_308_5_sva_dfm_1,
          sigmoid_table_309_5_sva_dfm_1, sigmoid_table_310_5_sva_dfm_1, sigmoid_table_311_5_sva_dfm_1,
          sigmoid_table_312_5_sva_dfm_1, sigmoid_table_313_5_sva_dfm_1, sigmoid_table_314_5_sva_dfm_1,
          sigmoid_table_315_5_sva_dfm_1, sigmoid_table_316_5_sva_dfm_1, sigmoid_table_317_5_sva_dfm_1,
          sigmoid_table_318_5_sva_dfm_1, sigmoid_table_319_5_sva_dfm_1, sigmoid_table_320_4_sva_dfm_1,
          sigmoid_table_321_4_sva_dfm_1, sigmoid_table_322_4_sva_dfm_1, sigmoid_table_323_4_sva_dfm_1,
          sigmoid_table_324_4_sva_dfm_1, sigmoid_table_325_4_sva_dfm_1, sigmoid_table_326_4_sva_dfm_1,
          sigmoid_table_327_4_sva_dfm_1, sigmoid_table_328_4_sva_dfm_1, sigmoid_table_329_4_sva_dfm_1,
          sigmoid_table_330_3_sva_dfm_1, sigmoid_table_331_3_sva_dfm_1, sigmoid_table_332_3_sva_dfm_1,
          sigmoid_table_333_3_sva_dfm_1, sigmoid_table_334_3_sva_dfm_1, sigmoid_table_335_2_sva_dfm_1,
          sigmoid_table_336_2_sva_dfm_1, sigmoid_table_337_1_sva_dfm_1, sigmoid_table_338_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_367_5_sva_dfm_1, sigmoid_table_368_5_sva_dfm_1,
          sigmoid_table_369_5_sva_dfm_1, sigmoid_table_370_5_sva_dfm_1, sigmoid_table_371_5_sva_dfm_1,
          sigmoid_table_372_5_sva_dfm_1, sigmoid_table_373_5_sva_dfm_1, sigmoid_table_374_5_sva_dfm_1,
          sigmoid_table_375_5_sva_dfm_1, sigmoid_table_376_5_sva_dfm_1, sigmoid_table_377_5_sva_dfm_1,
          sigmoid_table_378_4_sva_dfm_1, sigmoid_table_379_4_sva_dfm_1, sigmoid_table_380_4_sva_dfm_1,
          sigmoid_table_381_4_sva_dfm_1, sigmoid_table_382_4_sva_dfm_1, sigmoid_table_383_3_sva_dfm_1,
          sigmoid_table_384_3_sva_dfm_1, sigmoid_table_385_3_sva_dfm_1, sigmoid_table_386_2_sva_dfm_1,
          sigmoid_table_387_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_405_5_sva_dfm_1,
          sigmoid_table_406_5_sva_dfm_1, sigmoid_table_407_5_sva_dfm_1, sigmoid_table_408_5_sva_dfm_1,
          sigmoid_table_409_5_sva_dfm_1, sigmoid_table_410_5_sva_dfm_1, sigmoid_table_411_5_sva_dfm_1,
          sigmoid_table_412_4_sva_dfm_1, sigmoid_table_413_4_sva_dfm_1, sigmoid_table_414_4_sva_dfm_1,
          sigmoid_table_415_3_sva_dfm_1, sigmoid_table_416_3_sva_dfm_1, sigmoid_table_417_2_sva_dfm_1,
          sigmoid_table_418_0_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_431_5_sva_dfm_1, sigmoid_table_432_5_sva_dfm_1,
          sigmoid_table_433_5_sva_dfm_1, sigmoid_table_434_5_sva_dfm_1, sigmoid_table_435_5_sva_dfm_1,
          sigmoid_table_436_5_sva_dfm_1, sigmoid_table_437_4_sva_dfm_1, sigmoid_table_438_4_sva_dfm_1,
          sigmoid_table_439_3_sva_dfm_1, sigmoid_table_440_3_sva_dfm_1, sigmoid_table_441_2_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_452_5_sva_dfm_1,
          sigmoid_table_453_5_sva_dfm_1, sigmoid_table_454_5_sva_dfm_1, sigmoid_table_455_5_sva_dfm_1,
          sigmoid_table_456_5_sva_dfm_1, sigmoid_table_457_4_sva_dfm_1, sigmoid_table_458_4_sva_dfm_1,
          sigmoid_table_459_4_sva_dfm_1, sigmoid_table_460_3_sva_dfm_1, sigmoid_table_461_1_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_471_5_sva_dfm_1,
          sigmoid_table_472_5_sva_dfm_1, sigmoid_table_473_5_sva_dfm_1, sigmoid_table_474_5_sva_dfm_1,
          sigmoid_table_475_5_sva_dfm_1, sigmoid_table_476_4_sva_dfm_1, sigmoid_table_477_4_sva_dfm_1,
          sigmoid_table_478_3_sva_dfm_1, sigmoid_table_479_1_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_488_5_sva_dfm_1, sigmoid_table_489_5_sva_dfm_1,
          sigmoid_table_490_5_sva_dfm_1, sigmoid_table_491_5_sva_dfm_1, sigmoid_table_492_4_sva_dfm_1,
          sigmoid_table_493_4_sva_dfm_1, sigmoid_table_494_3_sva_dfm_1, sigmoid_table_495_2_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_504_5_sva_dfm_1,
          sigmoid_table_505_5_sva_dfm_1, sigmoid_table_506_5_sva_dfm_1, sigmoid_table_507_5_sva_dfm_1,
          sigmoid_table_508_4_sva_dfm_1, sigmoid_table_509_4_sva_dfm_1, sigmoid_table_510_3_sva_dfm_1,
          sigmoid_table_511_2_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_521_5_sva_dfm_1, sigmoid_table_522_5_sva_dfm_1,
          sigmoid_table_523_5_sva_dfm_1, sigmoid_table_524_5_sva_dfm_1, sigmoid_table_525_4_sva_dfm_1,
          sigmoid_table_526_4_sva_dfm_1, sigmoid_table_527_3_sva_dfm_1, sigmoid_table_528_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_537_5_sva_dfm_1,
          sigmoid_table_538_5_sva_dfm_1, sigmoid_table_539_5_sva_dfm_1, sigmoid_table_540_5_sva_dfm_1,
          sigmoid_table_541_4_sva_dfm_1, sigmoid_table_542_4_sva_dfm_1, sigmoid_table_543_3_sva_dfm_1,
          sigmoid_table_544_2_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, sigmoid_table_554_5_sva_dfm_1, sigmoid_table_555_5_sva_dfm_1,
          sigmoid_table_556_5_sva_dfm_1, sigmoid_table_557_5_sva_dfm_1, sigmoid_table_558_4_sva_dfm_1,
          sigmoid_table_559_4_sva_dfm_1, sigmoid_table_560_4_sva_dfm_1, sigmoid_table_561_3_sva_dfm_1,
          sigmoid_table_562_1_sva_dfm_1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, sigmoid_table_573_5_sva_dfm_1, sigmoid_table_574_5_sva_dfm_1,
          sigmoid_table_575_5_sva_dfm_1, sigmoid_table_576_5_sva_dfm_1, sigmoid_table_577_5_sva_dfm_1,
          sigmoid_table_578_4_sva_dfm_1, sigmoid_table_579_4_sva_dfm_1, sigmoid_table_580_3_sva_dfm_1,
          sigmoid_table_581_2_sva_dfm_1, sigmoid_table_582_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_594_5_sva_dfm_1,
          sigmoid_table_595_5_sva_dfm_1, sigmoid_table_596_5_sva_dfm_1, sigmoid_table_597_5_sva_dfm_1,
          sigmoid_table_598_5_sva_dfm_1, sigmoid_table_599_5_sva_dfm_1, sigmoid_table_600_4_sva_dfm_1,
          sigmoid_table_601_4_sva_dfm_1, sigmoid_table_602_4_sva_dfm_1, sigmoid_table_603_3_sva_dfm_1,
          sigmoid_table_604_3_sva_dfm_1, sigmoid_table_605_2_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          sigmoid_table_620_5_sva_dfm_1, sigmoid_table_621_5_sva_dfm_1, sigmoid_table_622_5_sva_dfm_1,
          sigmoid_table_623_5_sva_dfm_1, sigmoid_table_624_5_sva_dfm_1, sigmoid_table_625_5_sva_dfm_1,
          sigmoid_table_626_5_sva_dfm_1, sigmoid_table_627_5_sva_dfm_1, sigmoid_table_628_4_sva_dfm_1,
          sigmoid_table_629_4_sva_dfm_1, sigmoid_table_630_4_sva_dfm_1, sigmoid_table_631_4_sva_dfm_1,
          sigmoid_table_632_4_sva_dfm_1, sigmoid_table_633_3_sva_dfm_1, sigmoid_table_634_3_sva_dfm_1,
          sigmoid_table_635_2_sva_dfm_1, sigmoid_table_636_0_sva_dfm_1, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_658_5_sva_dfm_1,
          sigmoid_table_659_5_sva_dfm_1, sigmoid_table_660_5_sva_dfm_1, sigmoid_table_661_5_sva_dfm_1,
          sigmoid_table_662_5_sva_dfm_1, sigmoid_table_663_5_sva_dfm_1, sigmoid_table_664_5_sva_dfm_1,
          sigmoid_table_665_5_sva_dfm_1, sigmoid_table_666_5_sva_dfm_1, sigmoid_table_667_5_sva_dfm_1,
          sigmoid_table_668_5_sva_dfm_1, sigmoid_table_669_5_sva_dfm_1, sigmoid_table_670_4_sva_dfm_1,
          sigmoid_table_671_4_sva_dfm_1, sigmoid_table_672_4_sva_dfm_1, sigmoid_table_673_4_sva_dfm_1,
          sigmoid_table_674_4_sva_dfm_1, sigmoid_table_675_4_sva_dfm_1, sigmoid_table_676_4_sva_dfm_1,
          sigmoid_table_677_4_sva_dfm_1, sigmoid_table_678_3_sva_dfm_1, sigmoid_table_679_3_sva_dfm_1,
          sigmoid_table_680_3_sva_dfm_1, sigmoid_table_681_3_sva_dfm_1, sigmoid_table_682_2_sva_dfm_1,
          sigmoid_table_683_2_sva_dfm_1, sigmoid_table_684_1_sva_dfm_1, sigmoid_table_685_0_sva_dfm_1,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
          1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sigmoid_table_732_5_sva_dfm_1,
          sigmoid_table_733_5_sva_dfm_1, sigmoid_table_734_5_sva_dfm_1, sigmoid_table_735_5_sva_dfm_1,
          sigmoid_table_736_5_sva_dfm_1, sigmoid_table_737_5_sva_dfm_1, sigmoid_table_738_5_sva_dfm_1,
          sigmoid_table_739_5_sva_dfm_1, sigmoid_table_740_5_sva_dfm_1, sigmoid_table_741_5_sva_dfm_1,
          sigmoid_table_742_5_sva_dfm_1, sigmoid_table_743_5_sva_dfm_1, sigmoid_table_744_5_sva_dfm_1,
          sigmoid_table_745_5_sva_dfm_1, sigmoid_table_746_5_sva_dfm_1, sigmoid_table_747_5_sva_dfm_1,
          sigmoid_table_748_5_sva_dfm_1, sigmoid_table_749_5_sva_dfm_1, sigmoid_table_750_5_sva_dfm_1,
          sigmoid_table_751_5_sva_dfm_1, sigmoid_table_752_5_sva_dfm_1, sigmoid_table_753_5_sva_dfm_1,
          sigmoid_table_754_5_sva_dfm_1, sigmoid_table_755_5_sva_dfm_1, sigmoid_table_756_5_sva_dfm_1,
          sigmoid_table_757_5_sva_dfm_1, sigmoid_table_758_5_sva_dfm_1, sigmoid_table_759_5_sva_dfm_1,
          sigmoid_table_760_5_sva_dfm_1, sigmoid_table_761_5_sva_dfm_1, sigmoid_table_762_5_sva_dfm_1,
          sigmoid_table_763_5_sva_dfm_1, sigmoid_table_764_5_sva_dfm_1, sigmoid_table_765_5_sva_dfm_1,
          sigmoid_table_766_5_sva_dfm_1, sigmoid_table_767_5_sva_dfm_1, sigmoid_table_768_5_sva_dfm_1,
          sigmoid_table_769_5_sva_dfm_1, sigmoid_table_770_5_sva_dfm_1, sigmoid_table_771_5_sva_dfm_1,
          sigmoid_table_772_5_sva_dfm_1, sigmoid_table_773_5_sva_dfm_1, sigmoid_table_774_5_sva_dfm_1,
          sigmoid_table_775_5_sva_dfm_1, sigmoid_table_776_5_sva_dfm_1, sigmoid_table_777_5_sva_dfm_1,
          sigmoid_table_778_4_sva_dfm_1, sigmoid_table_779_4_sva_dfm_1, sigmoid_table_780_4_sva_dfm_1,
          sigmoid_table_781_4_sva_dfm_1, sigmoid_table_782_4_sva_dfm_1, sigmoid_table_783_4_sva_dfm_1,
          sigmoid_table_784_4_sva_dfm_1, sigmoid_table_785_4_sva_dfm_1, sigmoid_table_786_4_sva_dfm_1,
          sigmoid_table_787_4_sva_dfm_1, sigmoid_table_788_4_sva_dfm_1, sigmoid_table_789_4_sva_dfm_1,
          sigmoid_table_790_4_sva_dfm_1, sigmoid_table_791_4_sva_dfm_1, sigmoid_table_792_4_sva_dfm_1,
          sigmoid_table_793_4_sva_dfm_1, sigmoid_table_794_4_sva_dfm_1, sigmoid_table_795_4_sva_dfm_1,
          sigmoid_table_796_4_sva_dfm_1, sigmoid_table_797_4_sva_dfm_1, sigmoid_table_798_4_sva_dfm_1,
          sigmoid_table_799_4_sva_dfm_1, sigmoid_table_800_4_sva_dfm_1, sigmoid_table_801_4_sva_dfm_1,
          sigmoid_table_802_4_sva_dfm_1, sigmoid_table_803_4_sva_dfm_1, sigmoid_table_804_4_sva_dfm_1,
          sigmoid_table_805_4_sva_dfm_1, sigmoid_table_806_4_sva_dfm_1, sigmoid_table_807_4_sva_dfm_1,
          sigmoid_table_808_4_sva_dfm_1, sigmoid_table_809_4_sva_dfm_1, sigmoid_table_810_4_sva_dfm_1,
          sigmoid_table_811_4_sva_dfm_1, sigmoid_table_812_4_sva_dfm_1, sigmoid_table_813_4_sva_dfm_1,
          sigmoid_table_814_4_sva_dfm_1, sigmoid_table_815_4_sva_dfm_1, sigmoid_table_816_4_sva_dfm_1,
          sigmoid_table_817_4_sva_dfm_1, sigmoid_table_818_4_sva_dfm_1, sigmoid_table_819_4_sva_dfm_1,
          sigmoid_table_820_4_sva_dfm_1, sigmoid_table_821_4_sva_dfm_1, sigmoid_table_822_3_sva_dfm_1,
          sigmoid_table_823_3_sva_dfm_1, sigmoid_table_824_3_sva_dfm_1, sigmoid_table_825_3_sva_dfm_1,
          sigmoid_table_826_3_sva_dfm_1, sigmoid_table_827_3_sva_dfm_1, sigmoid_table_828_3_sva_dfm_1,
          sigmoid_table_829_3_sva_dfm_1, sigmoid_table_830_3_sva_dfm_1, sigmoid_table_831_3_sva_dfm_1,
          sigmoid_table_832_3_sva_dfm_1, sigmoid_table_833_3_sva_dfm_1, sigmoid_table_834_3_sva_dfm_1,
          sigmoid_table_835_3_sva_dfm_1, sigmoid_table_836_3_sva_dfm_1, sigmoid_table_837_3_sva_dfm_1,
          sigmoid_table_838_3_sva_dfm_1, sigmoid_table_839_3_sva_dfm_1, sigmoid_table_840_3_sva_dfm_1,
          sigmoid_table_841_3_sva_dfm_1, sigmoid_table_842_3_sva_dfm_1, sigmoid_table_843_3_sva_dfm_1,
          sigmoid_table_844_3_sva_dfm_1, sigmoid_table_845_3_sva_dfm_1, sigmoid_table_846_3_sva_dfm_1,
          sigmoid_table_847_3_sva_dfm_1, sigmoid_table_848_3_sva_dfm_1, sigmoid_table_849_3_sva_dfm_1,
          sigmoid_table_850_3_sva_dfm_1, sigmoid_table_851_3_sva_dfm_1, sigmoid_table_852_3_sva_dfm_1,
          sigmoid_table_853_3_sva_dfm_1, sigmoid_table_854_3_sva_dfm_1, sigmoid_table_855_3_sva_dfm_1,
          sigmoid_table_856_3_sva_dfm_1, sigmoid_table_857_3_sva_dfm_1, sigmoid_table_858_3_sva_dfm_1,
          sigmoid_table_859_3_sva_dfm_1, sigmoid_table_860_3_sva_dfm_1, sigmoid_table_861_3_sva_dfm_1,
          sigmoid_table_862_3_sva_dfm_1, sigmoid_table_863_3_sva_dfm_1, sigmoid_table_864_3_sva_dfm_1,
          sigmoid_table_865_3_sva_dfm_1, sigmoid_table_866_3_sva_dfm_1, sigmoid_table_867_2_sva_dfm_1,
          sigmoid_table_868_2_sva_dfm_1, sigmoid_table_869_2_sva_dfm_1, sigmoid_table_870_2_sva_dfm_1,
          sigmoid_table_871_2_sva_dfm_1, sigmoid_table_872_2_sva_dfm_1, sigmoid_table_873_2_sva_dfm_1,
          sigmoid_table_874_2_sva_dfm_1, sigmoid_table_875_2_sva_dfm_1, sigmoid_table_876_2_sva_dfm_1,
          sigmoid_table_877_2_sva_dfm_1, sigmoid_table_878_2_sva_dfm_1, sigmoid_table_879_2_sva_dfm_1,
          sigmoid_table_880_2_sva_dfm_1, sigmoid_table_881_2_sva_dfm_1, sigmoid_table_882_2_sva_dfm_1,
          sigmoid_table_883_2_sva_dfm_1, sigmoid_table_884_2_sva_dfm_1, sigmoid_table_885_2_sva_dfm_1,
          sigmoid_table_886_2_sva_dfm_1, sigmoid_table_887_2_sva_dfm_1, sigmoid_table_888_2_sva_dfm_1,
          sigmoid_table_889_2_sva_dfm_1, sigmoid_table_890_2_sva_dfm_1, sigmoid_table_891_2_sva_dfm_1,
          sigmoid_table_892_2_sva_dfm_1, sigmoid_table_893_2_sva_dfm_1, sigmoid_table_894_2_sva_dfm_1,
          sigmoid_table_895_2_sva_dfm_1, sigmoid_table_896_2_sva_dfm_1, sigmoid_table_897_2_sva_dfm_1,
          sigmoid_table_898_2_sva_dfm_1, sigmoid_table_899_2_sva_dfm_1, sigmoid_table_900_2_sva_dfm_1,
          sigmoid_table_901_2_sva_dfm_1, sigmoid_table_902_2_sva_dfm_1, sigmoid_table_903_2_sva_dfm_1,
          sigmoid_table_904_2_sva_dfm_1, sigmoid_table_905_2_sva_dfm_1, sigmoid_table_906_2_sva_dfm_1,
          sigmoid_table_907_2_sva_dfm_1, sigmoid_table_908_2_sva_dfm_1, sigmoid_table_909_2_sva_dfm_1,
          sigmoid_table_910_2_sva_dfm_1, sigmoid_table_911_1_sva_dfm_1, sigmoid_table_912_1_sva_dfm_1,
          sigmoid_table_913_1_sva_dfm_1, sigmoid_table_914_1_sva_dfm_1, sigmoid_table_915_1_sva_dfm_1,
          sigmoid_table_916_1_sva_dfm_1, sigmoid_table_917_1_sva_dfm_1, sigmoid_table_918_1_sva_dfm_1,
          sigmoid_table_919_1_sva_dfm_1, sigmoid_table_920_1_sva_dfm_1, sigmoid_table_921_1_sva_dfm_1,
          sigmoid_table_922_1_sva_dfm_1, sigmoid_table_923_1_sva_dfm_1, sigmoid_table_924_1_sva_dfm_1,
          sigmoid_table_925_1_sva_dfm_1, sigmoid_table_926_1_sva_dfm_1, sigmoid_table_927_1_sva_dfm_1,
          sigmoid_table_928_1_sva_dfm_1, sigmoid_table_929_1_sva_dfm_1, sigmoid_table_930_1_sva_dfm_1,
          sigmoid_table_931_1_sva_dfm_1, sigmoid_table_932_1_sva_dfm_1, sigmoid_table_933_1_sva_dfm_1,
          sigmoid_table_934_1_sva_dfm_1, sigmoid_table_935_1_sva_dfm_1, sigmoid_table_936_1_sva_dfm_1,
          sigmoid_table_937_1_sva_dfm_1, sigmoid_table_938_1_sva_dfm_1, sigmoid_table_939_1_sva_dfm_1,
          sigmoid_table_940_1_sva_dfm_1, sigmoid_table_941_1_sva_dfm_1, sigmoid_table_942_1_sva_dfm_1,
          sigmoid_table_943_1_sva_dfm_1, sigmoid_table_944_1_sva_dfm_1, sigmoid_table_945_1_sva_dfm_1,
          sigmoid_table_946_1_sva_dfm_1, sigmoid_table_947_1_sva_dfm_1, sigmoid_table_948_1_sva_dfm_1,
          sigmoid_table_949_1_sva_dfm_1, sigmoid_table_950_1_sva_dfm_1, sigmoid_table_951_1_sva_dfm_1,
          sigmoid_table_952_1_sva_dfm_1, sigmoid_table_953_1_sva_dfm_1, sigmoid_table_954_1_sva_dfm_1,
          sigmoid_table_955_0_sva_dfm_1, sigmoid_table_956_0_sva_dfm_1, sigmoid_table_957_0_sva_dfm_1,
          sigmoid_table_958_0_sva_dfm_1, sigmoid_table_959_0_sva_dfm_1, sigmoid_table_960_0_sva_dfm_1,
          sigmoid_table_961_0_sva_dfm_1, sigmoid_table_962_0_sva_dfm_1, sigmoid_table_963_0_sva_dfm_1,
          sigmoid_table_964_0_sva_dfm_1, sigmoid_table_965_0_sva_dfm_1, sigmoid_table_966_0_sva_dfm_1,
          sigmoid_table_967_0_sva_dfm_1, sigmoid_table_968_0_sva_dfm_1, sigmoid_table_969_0_sva_dfm_1,
          sigmoid_table_970_0_sva_dfm_1, sigmoid_table_971_0_sva_dfm_1, sigmoid_table_972_0_sva_dfm_1,
          sigmoid_table_973_0_sva_dfm_1, sigmoid_table_974_0_sva_dfm_1, sigmoid_table_975_0_sva_dfm_1,
          sigmoid_table_976_0_sva_dfm_1, sigmoid_table_977_0_sva_dfm_1, sigmoid_table_978_0_sva_dfm_1,
          sigmoid_table_979_0_sva_dfm_1, sigmoid_table_980_0_sva_dfm_1, sigmoid_table_981_0_sva_dfm_1,
          sigmoid_table_982_0_sva_dfm_1, sigmoid_table_983_0_sva_dfm_1, sigmoid_table_984_0_sva_dfm_1,
          sigmoid_table_985_0_sva_dfm_1, sigmoid_table_986_0_sva_dfm_1, sigmoid_table_987_0_sva_dfm_1,
          sigmoid_table_988_0_sva_dfm_1, sigmoid_table_989_0_sva_dfm_1, sigmoid_table_990_0_sva_dfm_1,
          sigmoid_table_991_0_sva_dfm_1, sigmoid_table_992_0_sva_dfm_1, sigmoid_table_993_0_sva_dfm_1,
          sigmoid_table_994_0_sva_dfm_1, sigmoid_table_995_0_sva_dfm_1, sigmoid_table_996_0_sva_dfm_1,
          sigmoid_table_997_0_sva_dfm_1, sigmoid_table_998_0_sva_dfm_1, sigmoid_table_999_0_sva_dfm_1,
          sigmoid_table_1000_0_sva_dfm_1, sigmoid_table_1001_0_sva_dfm_1, sigmoid_table_1002_0_sva_dfm_1,
          sigmoid_table_1003_0_sva_dfm_1, sigmoid_table_1004_0_sva_dfm_1, sigmoid_table_1005_0_sva_dfm_1,
          sigmoid_table_1006_0_sva_dfm_1, sigmoid_table_1007_0_sva_dfm_1, sigmoid_table_1008_0_sva_dfm_1,
          sigmoid_table_1009_0_sva_dfm_1, sigmoid_table_1010_0_sva_dfm_1, sigmoid_table_1011_0_sva_dfm_1,
          sigmoid_table_1012_0_sva_dfm_1, sigmoid_table_1013_0_sva_dfm_1, sigmoid_table_1014_0_sva_dfm_1,
          sigmoid_table_1015_0_sva_dfm_1, sigmoid_table_1016_0_sva_dfm_1, sigmoid_table_1017_0_sva_dfm_1,
          sigmoid_table_1018_0_sva_dfm_1, sigmoid_table_1019_0_sva_dfm_1, sigmoid_table_1020_0_sva_dfm_1,
          sigmoid_table_1021_0_sva_dfm_1, sigmoid_table_1022_0_sva_dfm_1, sigmoid_table_1023_0_sva_dfm_1,
          {for_for_or_1_itm , for_for_or_itm});
      initialized_sva <= initialized_sva | ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      sigmoid_table_1023_0_sva <= 1'b0;
      sigmoid_table_1022_0_sva <= 1'b0;
      sigmoid_table_1021_0_sva <= 1'b0;
      sigmoid_table_1020_0_sva <= 1'b0;
      sigmoid_table_1019_0_sva <= 1'b0;
      sigmoid_table_1018_0_sva <= 1'b0;
      sigmoid_table_1017_0_sva <= 1'b0;
      sigmoid_table_1016_0_sva <= 1'b0;
      sigmoid_table_1015_0_sva <= 1'b0;
      sigmoid_table_1014_0_sva <= 1'b0;
      sigmoid_table_1013_0_sva <= 1'b0;
      sigmoid_table_1012_0_sva <= 1'b0;
      sigmoid_table_1011_0_sva <= 1'b0;
      sigmoid_table_1010_0_sva <= 1'b0;
      sigmoid_table_1009_0_sva <= 1'b0;
      sigmoid_table_1008_0_sva <= 1'b0;
      sigmoid_table_1007_0_sva <= 1'b0;
      sigmoid_table_1006_0_sva <= 1'b0;
      sigmoid_table_1005_0_sva <= 1'b0;
      sigmoid_table_1004_0_sva <= 1'b0;
      sigmoid_table_1003_0_sva <= 1'b0;
      sigmoid_table_1002_0_sva <= 1'b0;
      sigmoid_table_1001_0_sva <= 1'b0;
      sigmoid_table_1000_0_sva <= 1'b0;
      sigmoid_table_999_0_sva <= 1'b0;
      sigmoid_table_998_0_sva <= 1'b0;
      sigmoid_table_997_0_sva <= 1'b0;
      sigmoid_table_996_0_sva <= 1'b0;
      sigmoid_table_995_0_sva <= 1'b0;
      sigmoid_table_994_0_sva <= 1'b0;
      sigmoid_table_993_0_sva <= 1'b0;
      sigmoid_table_992_0_sva <= 1'b0;
      sigmoid_table_991_0_sva <= 1'b0;
      sigmoid_table_990_0_sva <= 1'b0;
      sigmoid_table_989_0_sva <= 1'b0;
      sigmoid_table_988_0_sva <= 1'b0;
      sigmoid_table_987_0_sva <= 1'b0;
      sigmoid_table_986_0_sva <= 1'b0;
      sigmoid_table_985_0_sva <= 1'b0;
      sigmoid_table_984_0_sva <= 1'b0;
      sigmoid_table_983_0_sva <= 1'b0;
      sigmoid_table_982_0_sva <= 1'b0;
      sigmoid_table_981_0_sva <= 1'b0;
      sigmoid_table_980_0_sva <= 1'b0;
      sigmoid_table_979_0_sva <= 1'b0;
      sigmoid_table_978_0_sva <= 1'b0;
      sigmoid_table_977_0_sva <= 1'b0;
      sigmoid_table_976_0_sva <= 1'b0;
      sigmoid_table_975_0_sva <= 1'b0;
      sigmoid_table_974_0_sva <= 1'b0;
      sigmoid_table_973_0_sva <= 1'b0;
      sigmoid_table_972_0_sva <= 1'b0;
      sigmoid_table_971_0_sva <= 1'b0;
      sigmoid_table_970_0_sva <= 1'b0;
      sigmoid_table_969_0_sva <= 1'b0;
      sigmoid_table_968_0_sva <= 1'b0;
      sigmoid_table_967_0_sva <= 1'b0;
      sigmoid_table_966_0_sva <= 1'b0;
      sigmoid_table_965_0_sva <= 1'b0;
      sigmoid_table_964_0_sva <= 1'b0;
      sigmoid_table_963_0_sva <= 1'b0;
      sigmoid_table_962_0_sva <= 1'b0;
      sigmoid_table_961_0_sva <= 1'b0;
      sigmoid_table_960_0_sva <= 1'b0;
      sigmoid_table_959_0_sva <= 1'b0;
      sigmoid_table_958_0_sva <= 1'b0;
      sigmoid_table_957_0_sva <= 1'b0;
      sigmoid_table_956_0_sva <= 1'b0;
      sigmoid_table_955_0_sva <= 1'b0;
      sigmoid_table_954_1_sva <= 1'b0;
      sigmoid_table_953_1_sva <= 1'b0;
      sigmoid_table_952_1_sva <= 1'b0;
      sigmoid_table_951_1_sva <= 1'b0;
      sigmoid_table_950_1_sva <= 1'b0;
      sigmoid_table_949_1_sva <= 1'b0;
      sigmoid_table_948_1_sva <= 1'b0;
      sigmoid_table_947_1_sva <= 1'b0;
      sigmoid_table_946_1_sva <= 1'b0;
      sigmoid_table_945_1_sva <= 1'b0;
      sigmoid_table_944_1_sva <= 1'b0;
      sigmoid_table_943_1_sva <= 1'b0;
      sigmoid_table_942_1_sva <= 1'b0;
      sigmoid_table_941_1_sva <= 1'b0;
      sigmoid_table_940_1_sva <= 1'b0;
      sigmoid_table_939_1_sva <= 1'b0;
      sigmoid_table_938_1_sva <= 1'b0;
      sigmoid_table_937_1_sva <= 1'b0;
      sigmoid_table_936_1_sva <= 1'b0;
      sigmoid_table_935_1_sva <= 1'b0;
      sigmoid_table_934_1_sva <= 1'b0;
      sigmoid_table_933_1_sva <= 1'b0;
      sigmoid_table_932_1_sva <= 1'b0;
      sigmoid_table_931_1_sva <= 1'b0;
      sigmoid_table_930_1_sva <= 1'b0;
      sigmoid_table_929_1_sva <= 1'b0;
      sigmoid_table_928_1_sva <= 1'b0;
      sigmoid_table_927_1_sva <= 1'b0;
      sigmoid_table_926_1_sva <= 1'b0;
      sigmoid_table_925_1_sva <= 1'b0;
      sigmoid_table_924_1_sva <= 1'b0;
      sigmoid_table_923_1_sva <= 1'b0;
      sigmoid_table_922_1_sva <= 1'b0;
      sigmoid_table_921_1_sva <= 1'b0;
      sigmoid_table_920_1_sva <= 1'b0;
      sigmoid_table_919_1_sva <= 1'b0;
      sigmoid_table_918_1_sva <= 1'b0;
      sigmoid_table_917_1_sva <= 1'b0;
      sigmoid_table_916_1_sva <= 1'b0;
      sigmoid_table_915_1_sva <= 1'b0;
      sigmoid_table_914_1_sva <= 1'b0;
      sigmoid_table_913_1_sva <= 1'b0;
      sigmoid_table_912_1_sva <= 1'b0;
      sigmoid_table_911_1_sva <= 1'b0;
      sigmoid_table_910_2_sva <= 1'b0;
      sigmoid_table_909_2_sva <= 1'b0;
      sigmoid_table_908_2_sva <= 1'b0;
      sigmoid_table_907_2_sva <= 1'b0;
      sigmoid_table_906_2_sva <= 1'b0;
      sigmoid_table_905_2_sva <= 1'b0;
      sigmoid_table_904_2_sva <= 1'b0;
      sigmoid_table_903_2_sva <= 1'b0;
      sigmoid_table_902_2_sva <= 1'b0;
      sigmoid_table_901_2_sva <= 1'b0;
      sigmoid_table_900_2_sva <= 1'b0;
      sigmoid_table_899_2_sva <= 1'b0;
      sigmoid_table_898_2_sva <= 1'b0;
      sigmoid_table_897_2_sva <= 1'b0;
      sigmoid_table_896_2_sva <= 1'b0;
      sigmoid_table_895_2_sva <= 1'b0;
      sigmoid_table_894_2_sva <= 1'b0;
      sigmoid_table_893_2_sva <= 1'b0;
      sigmoid_table_892_2_sva <= 1'b0;
      sigmoid_table_891_2_sva <= 1'b0;
      sigmoid_table_890_2_sva <= 1'b0;
      sigmoid_table_889_2_sva <= 1'b0;
      sigmoid_table_888_2_sva <= 1'b0;
      sigmoid_table_887_2_sva <= 1'b0;
      sigmoid_table_886_2_sva <= 1'b0;
      sigmoid_table_885_2_sva <= 1'b0;
      sigmoid_table_884_2_sva <= 1'b0;
      sigmoid_table_883_2_sva <= 1'b0;
      sigmoid_table_882_2_sva <= 1'b0;
      sigmoid_table_881_2_sva <= 1'b0;
      sigmoid_table_880_2_sva <= 1'b0;
      sigmoid_table_879_2_sva <= 1'b0;
      sigmoid_table_878_2_sva <= 1'b0;
      sigmoid_table_877_2_sva <= 1'b0;
      sigmoid_table_876_2_sva <= 1'b0;
      sigmoid_table_875_2_sva <= 1'b0;
      sigmoid_table_874_2_sva <= 1'b0;
      sigmoid_table_873_2_sva <= 1'b0;
      sigmoid_table_872_2_sva <= 1'b0;
      sigmoid_table_871_2_sva <= 1'b0;
      sigmoid_table_870_2_sva <= 1'b0;
      sigmoid_table_869_2_sva <= 1'b0;
      sigmoid_table_868_2_sva <= 1'b0;
      sigmoid_table_867_2_sva <= 1'b0;
      sigmoid_table_866_0_sva <= 1'b0;
      sigmoid_table_866_3_sva <= 1'b0;
      sigmoid_table_865_0_sva <= 1'b0;
      sigmoid_table_865_3_sva <= 1'b0;
      sigmoid_table_864_0_sva <= 1'b0;
      sigmoid_table_864_3_sva <= 1'b0;
      sigmoid_table_863_0_sva <= 1'b0;
      sigmoid_table_863_3_sva <= 1'b0;
      sigmoid_table_862_0_sva <= 1'b0;
      sigmoid_table_862_3_sva <= 1'b0;
      sigmoid_table_861_0_sva <= 1'b0;
      sigmoid_table_861_3_sva <= 1'b0;
      sigmoid_table_860_0_sva <= 1'b0;
      sigmoid_table_860_3_sva <= 1'b0;
      sigmoid_table_859_0_sva <= 1'b0;
      sigmoid_table_859_3_sva <= 1'b0;
      sigmoid_table_858_0_sva <= 1'b0;
      sigmoid_table_858_3_sva <= 1'b0;
      sigmoid_table_857_0_sva <= 1'b0;
      sigmoid_table_857_3_sva <= 1'b0;
      sigmoid_table_856_0_sva <= 1'b0;
      sigmoid_table_856_3_sva <= 1'b0;
      sigmoid_table_855_0_sva <= 1'b0;
      sigmoid_table_855_3_sva <= 1'b0;
      sigmoid_table_854_0_sva <= 1'b0;
      sigmoid_table_854_3_sva <= 1'b0;
      sigmoid_table_853_0_sva <= 1'b0;
      sigmoid_table_853_3_sva <= 1'b0;
      sigmoid_table_852_3_sva <= 1'b0;
      sigmoid_table_851_3_sva <= 1'b0;
      sigmoid_table_850_3_sva <= 1'b0;
      sigmoid_table_849_3_sva <= 1'b0;
      sigmoid_table_848_3_sva <= 1'b0;
      sigmoid_table_847_3_sva <= 1'b0;
      sigmoid_table_846_3_sva <= 1'b0;
      sigmoid_table_845_3_sva <= 1'b0;
      sigmoid_table_844_3_sva <= 1'b0;
      sigmoid_table_843_3_sva <= 1'b0;
      sigmoid_table_842_3_sva <= 1'b0;
      sigmoid_table_841_3_sva <= 1'b0;
      sigmoid_table_840_3_sva <= 1'b0;
      sigmoid_table_839_3_sva <= 1'b0;
      sigmoid_table_838_3_sva <= 1'b0;
      sigmoid_table_837_3_sva <= 1'b0;
      sigmoid_table_836_3_sva <= 1'b0;
      sigmoid_table_835_3_sva <= 1'b0;
      sigmoid_table_834_3_sva <= 1'b0;
      sigmoid_table_833_3_sva <= 1'b0;
      sigmoid_table_832_3_sva <= 1'b0;
      sigmoid_table_831_3_sva <= 1'b0;
      sigmoid_table_830_3_sva <= 1'b0;
      sigmoid_table_829_3_sva <= 1'b0;
      sigmoid_table_828_3_sva <= 1'b0;
      sigmoid_table_827_3_sva <= 1'b0;
      sigmoid_table_826_3_sva <= 1'b0;
      sigmoid_table_825_3_sva <= 1'b0;
      sigmoid_table_824_3_sva <= 1'b0;
      sigmoid_table_823_3_sva <= 1'b0;
      sigmoid_table_822_3_sva <= 1'b0;
      sigmoid_table_821_0_sva <= 1'b0;
      sigmoid_table_821_4_sva <= 1'b0;
      sigmoid_table_820_0_sva <= 1'b0;
      sigmoid_table_820_4_sva <= 1'b0;
      sigmoid_table_819_0_sva <= 1'b0;
      sigmoid_table_819_4_sva <= 1'b0;
      sigmoid_table_818_0_sva <= 1'b0;
      sigmoid_table_818_4_sva <= 1'b0;
      sigmoid_table_817_0_sva <= 1'b0;
      sigmoid_table_817_4_sva <= 1'b0;
      sigmoid_table_816_0_sva <= 1'b0;
      sigmoid_table_816_4_sva <= 1'b0;
      sigmoid_table_815_0_sva <= 1'b0;
      sigmoid_table_815_4_sva <= 1'b0;
      sigmoid_table_814_1_sva <= 1'b0;
      sigmoid_table_814_4_sva <= 1'b0;
      sigmoid_table_813_1_sva <= 1'b0;
      sigmoid_table_813_4_sva <= 1'b0;
      sigmoid_table_812_1_sva <= 1'b0;
      sigmoid_table_812_4_sva <= 1'b0;
      sigmoid_table_811_1_sva <= 1'b0;
      sigmoid_table_811_4_sva <= 1'b0;
      sigmoid_table_810_1_sva <= 1'b0;
      sigmoid_table_810_4_sva <= 1'b0;
      sigmoid_table_809_1_sva <= 1'b0;
      sigmoid_table_809_4_sva <= 1'b0;
      sigmoid_table_808_1_sva <= 1'b0;
      sigmoid_table_808_4_sva <= 1'b0;
      sigmoid_table_807_4_sva <= 1'b0;
      sigmoid_table_806_4_sva <= 1'b0;
      sigmoid_table_805_4_sva <= 1'b0;
      sigmoid_table_804_4_sva <= 1'b0;
      sigmoid_table_803_4_sva <= 1'b0;
      sigmoid_table_802_4_sva <= 1'b0;
      sigmoid_table_801_4_sva <= 1'b0;
      sigmoid_table_800_4_sva <= 1'b0;
      sigmoid_table_799_4_sva <= 1'b0;
      sigmoid_table_798_4_sva <= 1'b0;
      sigmoid_table_797_4_sva <= 1'b0;
      sigmoid_table_796_4_sva <= 1'b0;
      sigmoid_table_795_0_sva <= 1'b0;
      sigmoid_table_795_4_sva <= 1'b0;
      sigmoid_table_794_0_sva <= 1'b0;
      sigmoid_table_794_4_sva <= 1'b0;
      sigmoid_table_793_0_sva <= 1'b0;
      sigmoid_table_793_4_sva <= 1'b0;
      sigmoid_table_792_0_sva <= 1'b0;
      sigmoid_table_792_4_sva <= 1'b0;
      sigmoid_table_791_0_sva <= 1'b0;
      sigmoid_table_791_4_sva <= 1'b0;
      sigmoid_table_790_4_sva <= 1'b0;
      sigmoid_table_789_4_sva <= 1'b0;
      sigmoid_table_788_4_sva <= 1'b0;
      sigmoid_table_787_4_sva <= 1'b0;
      sigmoid_table_786_4_sva <= 1'b0;
      sigmoid_table_785_4_sva <= 1'b0;
      sigmoid_table_784_4_sva <= 1'b0;
      sigmoid_table_783_4_sva <= 1'b0;
      sigmoid_table_782_4_sva <= 1'b0;
      sigmoid_table_781_4_sva <= 1'b0;
      sigmoid_table_780_4_sva <= 1'b0;
      sigmoid_table_779_4_sva <= 1'b0;
      sigmoid_table_778_4_sva <= 1'b0;
      sigmoid_table_777_0_sva <= 1'b0;
      sigmoid_table_777_5_sva <= 1'b0;
      sigmoid_table_776_0_sva <= 1'b0;
      sigmoid_table_776_5_sva <= 1'b0;
      sigmoid_table_775_0_sva <= 1'b0;
      sigmoid_table_775_5_sva <= 1'b0;
      sigmoid_table_774_0_sva <= 1'b0;
      sigmoid_table_774_5_sva <= 1'b0;
      sigmoid_table_773_1_sva <= 1'b0;
      sigmoid_table_773_5_sva <= 1'b0;
      sigmoid_table_772_1_sva <= 1'b0;
      sigmoid_table_772_5_sva <= 1'b0;
      sigmoid_table_771_1_sva <= 1'b0;
      sigmoid_table_771_5_sva <= 1'b0;
      sigmoid_table_770_1_sva <= 1'b0;
      sigmoid_table_770_5_sva <= 1'b0;
      sigmoid_table_769_2_sva <= 1'b0;
      sigmoid_table_769_5_sva <= 1'b0;
      sigmoid_table_768_2_sva <= 1'b0;
      sigmoid_table_768_5_sva <= 1'b0;
      sigmoid_table_767_2_sva <= 1'b0;
      sigmoid_table_767_5_sva <= 1'b0;
      sigmoid_table_766_2_sva <= 1'b0;
      sigmoid_table_766_5_sva <= 1'b0;
      sigmoid_table_765_2_sva <= 1'b0;
      sigmoid_table_765_5_sva <= 1'b0;
      sigmoid_table_764_2_sva <= 1'b0;
      sigmoid_table_764_5_sva <= 1'b0;
      sigmoid_table_763_2_sva <= 1'b0;
      sigmoid_table_763_5_sva <= 1'b0;
      sigmoid_table_762_0_sva <= 1'b0;
      sigmoid_table_762_5_sva <= 1'b0;
      sigmoid_table_761_0_sva <= 1'b0;
      sigmoid_table_761_5_sva <= 1'b0;
      sigmoid_table_760_0_sva <= 1'b0;
      sigmoid_table_760_5_sva <= 1'b0;
      sigmoid_table_759_5_sva <= 1'b0;
      sigmoid_table_758_5_sva <= 1'b0;
      sigmoid_table_757_5_sva <= 1'b0;
      sigmoid_table_756_5_sva <= 1'b0;
      sigmoid_table_755_5_sva <= 1'b0;
      sigmoid_table_754_5_sva <= 1'b0;
      sigmoid_table_753_5_sva <= 1'b0;
      sigmoid_table_752_5_sva <= 1'b0;
      sigmoid_table_751_5_sva <= 1'b0;
      sigmoid_table_750_0_sva <= 1'b0;
      sigmoid_table_750_5_sva <= 1'b0;
      sigmoid_table_749_0_sva <= 1'b0;
      sigmoid_table_749_5_sva <= 1'b0;
      sigmoid_table_748_0_sva <= 1'b0;
      sigmoid_table_748_5_sva <= 1'b0;
      sigmoid_table_747_1_sva <= 1'b0;
      sigmoid_table_747_5_sva <= 1'b0;
      sigmoid_table_746_1_sva <= 1'b0;
      sigmoid_table_746_5_sva <= 1'b0;
      sigmoid_table_745_5_sva <= 1'b0;
      sigmoid_table_744_5_sva <= 1'b0;
      sigmoid_table_743_5_sva <= 1'b0;
      sigmoid_table_742_5_sva <= 1'b0;
      sigmoid_table_741_5_sva <= 1'b0;
      sigmoid_table_740_0_sva <= 1'b0;
      sigmoid_table_740_5_sva <= 1'b0;
      sigmoid_table_739_0_sva <= 1'b0;
      sigmoid_table_739_5_sva <= 1'b0;
      sigmoid_table_738_5_sva <= 1'b0;
      sigmoid_table_737_5_sva <= 1'b0;
      sigmoid_table_736_5_sva <= 1'b0;
      sigmoid_table_735_5_sva <= 1'b0;
      sigmoid_table_734_5_sva <= 1'b0;
      sigmoid_table_733_5_sva <= 1'b0;
      sigmoid_table_732_5_sva <= 1'b0;
      sigmoid_table_731_0_sva <= 1'b0;
      sigmoid_table_731_6_sva <= 1'b0;
      sigmoid_table_730_0_sva <= 1'b0;
      sigmoid_table_730_6_sva <= 1'b0;
      sigmoid_table_729_1_sva <= 1'b0;
      sigmoid_table_729_6_sva <= 1'b0;
      sigmoid_table_728_1_sva <= 1'b0;
      sigmoid_table_728_6_sva <= 1'b0;
      sigmoid_table_727_2_sva <= 1'b0;
      sigmoid_table_727_6_sva <= 1'b0;
      sigmoid_table_726_2_sva <= 1'b0;
      sigmoid_table_726_6_sva <= 1'b0;
      sigmoid_table_725_2_sva <= 1'b0;
      sigmoid_table_725_6_sva <= 1'b0;
      sigmoid_table_724_2_sva <= 1'b0;
      sigmoid_table_724_6_sva <= 1'b0;
      sigmoid_table_723_0_sva <= 1'b0;
      sigmoid_table_723_3_sva <= 1'b0;
      sigmoid_table_723_6_sva <= 1'b0;
      sigmoid_table_722_3_sva <= 1'b0;
      sigmoid_table_722_6_sva <= 1'b0;
      sigmoid_table_721_3_sva <= 1'b0;
      sigmoid_table_721_6_sva <= 1'b0;
      sigmoid_table_720_3_sva <= 1'b0;
      sigmoid_table_720_6_sva <= 1'b0;
      sigmoid_table_719_3_sva <= 1'b0;
      sigmoid_table_719_6_sva <= 1'b0;
      sigmoid_table_718_3_sva <= 1'b0;
      sigmoid_table_718_6_sva <= 1'b0;
      sigmoid_table_717_3_sva <= 1'b0;
      sigmoid_table_717_6_sva <= 1'b0;
      sigmoid_table_716_0_sva <= 1'b0;
      sigmoid_table_716_6_sva <= 1'b0;
      sigmoid_table_715_1_sva <= 1'b0;
      sigmoid_table_715_6_sva <= 1'b0;
      sigmoid_table_714_1_sva <= 1'b0;
      sigmoid_table_714_6_sva <= 1'b0;
      sigmoid_table_713_6_sva <= 1'b0;
      sigmoid_table_712_6_sva <= 1'b0;
      sigmoid_table_711_6_sva <= 1'b0;
      sigmoid_table_710_0_sva <= 1'b0;
      sigmoid_table_710_6_sva <= 1'b0;
      sigmoid_table_709_6_sva <= 1'b0;
      sigmoid_table_708_6_sva <= 1'b0;
      sigmoid_table_707_6_sva <= 1'b0;
      sigmoid_table_706_6_sva <= 1'b0;
      sigmoid_table_705_6_sva <= 1'b0;
      sigmoid_table_704_0_sva <= 1'b0;
      sigmoid_table_704_6_sva <= 1'b0;
      sigmoid_table_703_1_sva <= 1'b0;
      sigmoid_table_703_6_sva <= 1'b0;
      sigmoid_table_702_2_sva <= 1'b0;
      sigmoid_table_702_6_sva <= 1'b0;
      sigmoid_table_701_2_sva <= 1'b0;
      sigmoid_table_701_6_sva <= 1'b0;
      sigmoid_table_700_2_sva <= 1'b0;
      sigmoid_table_700_6_sva <= 1'b0;
      sigmoid_table_699_0_sva <= 1'b0;
      sigmoid_table_699_6_sva <= 1'b0;
      sigmoid_table_698_6_sva <= 1'b0;
      sigmoid_table_697_6_sva <= 1'b0;
      sigmoid_table_696_6_sva <= 1'b0;
      sigmoid_table_695_6_sva <= 1'b0;
      sigmoid_table_694_0_sva <= 1'b0;
      sigmoid_table_694_6_sva <= 1'b0;
      sigmoid_table_693_1_sva <= 1'b0;
      sigmoid_table_693_6_sva <= 1'b0;
      sigmoid_table_692_6_sva <= 1'b0;
      sigmoid_table_691_6_sva <= 1'b0;
      sigmoid_table_690_6_sva <= 1'b0;
      sigmoid_table_689_0_sva <= 1'b0;
      sigmoid_table_689_6_sva <= 1'b0;
      sigmoid_table_688_6_sva <= 1'b0;
      sigmoid_table_687_6_sva <= 1'b0;
      sigmoid_table_686_6_sva <= 1'b0;
      sigmoid_table_685_0_sva <= 1'b0;
      sigmoid_table_685_7_sva <= 1'b0;
      sigmoid_table_684_1_sva <= 1'b0;
      sigmoid_table_684_7_sva <= 1'b0;
      sigmoid_table_683_2_sva <= 1'b0;
      sigmoid_table_683_7_sva <= 1'b0;
      sigmoid_table_682_2_sva <= 1'b0;
      sigmoid_table_682_7_sva <= 1'b0;
      sigmoid_table_681_0_sva <= 1'b0;
      sigmoid_table_681_3_sva <= 1'b0;
      sigmoid_table_681_7_sva <= 1'b0;
      sigmoid_table_680_3_sva <= 1'b0;
      sigmoid_table_680_7_sva <= 1'b0;
      sigmoid_table_679_3_sva <= 1'b0;
      sigmoid_table_679_7_sva <= 1'b0;
      sigmoid_table_678_3_sva <= 1'b0;
      sigmoid_table_678_7_sva <= 1'b0;
      sigmoid_table_677_0_sva <= 1'b0;
      sigmoid_table_677_4_sva <= 1'b0;
      sigmoid_table_677_7_sva <= 1'b0;
      sigmoid_table_676_1_sva <= 1'b0;
      sigmoid_table_676_4_sva <= 1'b0;
      sigmoid_table_676_7_sva <= 1'b0;
      sigmoid_table_675_4_sva <= 1'b0;
      sigmoid_table_675_7_sva <= 1'b0;
      sigmoid_table_674_4_sva <= 1'b0;
      sigmoid_table_674_7_sva <= 1'b0;
      sigmoid_table_673_0_sva <= 1'b0;
      sigmoid_table_673_4_sva <= 1'b0;
      sigmoid_table_673_7_sva <= 1'b0;
      sigmoid_table_672_4_sva <= 1'b0;
      sigmoid_table_672_7_sva <= 1'b0;
      sigmoid_table_671_4_sva <= 1'b0;
      sigmoid_table_671_7_sva <= 1'b0;
      sigmoid_table_670_4_sva <= 1'b0;
      sigmoid_table_670_7_sva <= 1'b0;
      sigmoid_table_669_1_sva <= 1'b0;
      sigmoid_table_669_7_sva <= 1'b0;
      sigmoid_table_668_2_sva <= 1'b0;
      sigmoid_table_668_7_sva <= 1'b0;
      sigmoid_table_667_2_sva <= 1'b0;
      sigmoid_table_667_7_sva <= 1'b0;
      sigmoid_table_666_0_sva <= 1'b0;
      sigmoid_table_666_7_sva <= 1'b0;
      sigmoid_table_665_7_sva <= 1'b0;
      sigmoid_table_664_7_sva <= 1'b0;
      sigmoid_table_663_0_sva <= 1'b0;
      sigmoid_table_663_7_sva <= 1'b0;
      sigmoid_table_662_1_sva <= 1'b0;
      sigmoid_table_662_7_sva <= 1'b0;
      sigmoid_table_661_7_sva <= 1'b0;
      sigmoid_table_660_0_sva <= 1'b0;
      sigmoid_table_660_7_sva <= 1'b0;
      sigmoid_table_659_7_sva <= 1'b0;
      sigmoid_table_658_7_sva <= 1'b0;
      sigmoid_table_657_0_sva <= 1'b0;
      sigmoid_table_657_7_sva <= 1'b0;
      sigmoid_table_656_1_sva <= 1'b0;
      sigmoid_table_656_7_sva <= 1'b0;
      sigmoid_table_655_2_sva <= 1'b0;
      sigmoid_table_655_7_sva <= 1'b0;
      sigmoid_table_654_0_sva <= 1'b0;
      sigmoid_table_654_3_sva <= 1'b0;
      sigmoid_table_654_7_sva <= 1'b0;
      sigmoid_table_653_3_sva <= 1'b0;
      sigmoid_table_653_7_sva <= 1'b0;
      sigmoid_table_652_3_sva <= 1'b0;
      sigmoid_table_652_7_sva <= 1'b0;
      sigmoid_table_651_0_sva <= 1'b0;
      sigmoid_table_651_7_sva <= 1'b0;
      sigmoid_table_650_7_sva <= 1'b0;
      sigmoid_table_649_7_sva <= 1'b0;
      sigmoid_table_648_7_sva <= 1'b0;
      sigmoid_table_647_7_sva <= 1'b0;
      sigmoid_table_646_0_sva <= 1'b0;
      sigmoid_table_646_7_sva <= 1'b0;
      sigmoid_table_645_1_sva <= 1'b0;
      sigmoid_table_645_7_sva <= 1'b0;
      sigmoid_table_644_2_sva <= 1'b0;
      sigmoid_table_644_7_sva <= 1'b0;
      sigmoid_table_643_7_sva <= 1'b0;
      sigmoid_table_642_7_sva <= 1'b0;
      sigmoid_table_641_0_sva <= 1'b0;
      sigmoid_table_641_7_sva <= 1'b0;
      sigmoid_table_640_7_sva <= 1'b0;
      sigmoid_table_639_7_sva <= 1'b0;
      sigmoid_table_638_7_sva <= 1'b0;
      sigmoid_table_637_7_sva <= 1'b0;
      sigmoid_table_636_0_sva <= 1'b0;
      sigmoid_table_636_8_sva <= 1'b0;
      sigmoid_table_635_2_sva <= 1'b0;
      sigmoid_table_635_8_sva <= 1'b0;
      sigmoid_table_634_0_sva <= 1'b0;
      sigmoid_table_634_3_sva <= 1'b0;
      sigmoid_table_634_8_sva <= 1'b0;
      sigmoid_table_633_3_sva <= 1'b0;
      sigmoid_table_633_8_sva <= 1'b0;
      sigmoid_table_632_0_sva <= 1'b0;
      sigmoid_table_632_4_sva <= 1'b0;
      sigmoid_table_632_8_sva <= 1'b0;
      sigmoid_table_631_4_sva <= 1'b0;
      sigmoid_table_631_8_sva <= 1'b0;
      sigmoid_table_630_4_sva <= 1'b0;
      sigmoid_table_630_8_sva <= 1'b0;
      sigmoid_table_629_4_sva <= 1'b0;
      sigmoid_table_629_8_sva <= 1'b0;
      sigmoid_table_628_4_sva <= 1'b0;
      sigmoid_table_628_8_sva <= 1'b0;
      sigmoid_table_627_1_sva <= 1'b0;
      sigmoid_table_627_5_sva <= 1'b0;
      sigmoid_table_627_8_sva <= 1'b0;
      sigmoid_table_626_2_sva <= 1'b0;
      sigmoid_table_626_5_sva <= 1'b0;
      sigmoid_table_626_8_sva <= 1'b0;
      sigmoid_table_625_5_sva <= 1'b0;
      sigmoid_table_625_8_sva <= 1'b0;
      sigmoid_table_624_5_sva <= 1'b0;
      sigmoid_table_624_8_sva <= 1'b0;
      sigmoid_table_623_1_sva <= 1'b0;
      sigmoid_table_623_5_sva <= 1'b0;
      sigmoid_table_623_8_sva <= 1'b0;
      sigmoid_table_622_5_sva <= 1'b0;
      sigmoid_table_622_8_sva <= 1'b0;
      sigmoid_table_621_5_sva <= 1'b0;
      sigmoid_table_621_8_sva <= 1'b0;
      sigmoid_table_620_5_sva <= 1'b0;
      sigmoid_table_620_8_sva <= 1'b0;
      sigmoid_table_619_1_sva <= 1'b0;
      sigmoid_table_619_8_sva <= 1'b0;
      sigmoid_table_618_0_sva <= 1'b0;
      sigmoid_table_618_3_sva <= 1'b0;
      sigmoid_table_618_8_sva <= 1'b0;
      sigmoid_table_617_3_sva <= 1'b0;
      sigmoid_table_617_8_sva <= 1'b0;
      sigmoid_table_616_0_sva <= 1'b0;
      sigmoid_table_616_8_sva <= 1'b0;
      sigmoid_table_615_8_sva <= 1'b0;
      sigmoid_table_614_0_sva <= 1'b0;
      sigmoid_table_614_8_sva <= 1'b0;
      sigmoid_table_613_8_sva <= 1'b0;
      sigmoid_table_612_1_sva <= 1'b0;
      sigmoid_table_612_8_sva <= 1'b0;
      sigmoid_table_611_2_sva <= 1'b0;
      sigmoid_table_611_8_sva <= 1'b0;
      sigmoid_table_610_8_sva <= 1'b0;
      sigmoid_table_609_0_sva <= 1'b0;
      sigmoid_table_609_8_sva <= 1'b0;
      sigmoid_table_608_8_sva <= 1'b0;
      sigmoid_table_607_8_sva <= 1'b0;
      sigmoid_table_606_8_sva <= 1'b0;
      sigmoid_table_605_2_sva <= 1'b0;
      sigmoid_table_605_8_sva <= 1'b0;
      sigmoid_table_604_0_sva <= 1'b0;
      sigmoid_table_604_3_sva <= 1'b0;
      sigmoid_table_604_8_sva <= 1'b0;
      sigmoid_table_603_3_sva <= 1'b0;
      sigmoid_table_603_8_sva <= 1'b0;
      sigmoid_table_602_1_sva <= 1'b0;
      sigmoid_table_602_4_sva <= 1'b0;
      sigmoid_table_602_8_sva <= 1'b0;
      sigmoid_table_601_0_sva <= 1'b0;
      sigmoid_table_601_4_sva <= 1'b0;
      sigmoid_table_601_8_sva <= 1'b0;
      sigmoid_table_600_4_sva <= 1'b0;
      sigmoid_table_600_8_sva <= 1'b0;
      sigmoid_table_599_1_sva <= 1'b0;
      sigmoid_table_599_8_sva <= 1'b0;
      sigmoid_table_598_2_sva <= 1'b0;
      sigmoid_table_598_8_sva <= 1'b0;
      sigmoid_table_597_8_sva <= 1'b0;
      sigmoid_table_596_1_sva <= 1'b0;
      sigmoid_table_596_8_sva <= 1'b0;
      sigmoid_table_595_8_sva <= 1'b0;
      sigmoid_table_594_8_sva <= 1'b0;
      sigmoid_table_593_1_sva <= 1'b0;
      sigmoid_table_593_8_sva <= 1'b0;
      sigmoid_table_592_0_sva <= 1'b0;
      sigmoid_table_592_3_sva <= 1'b0;
      sigmoid_table_592_8_sva <= 1'b0;
      sigmoid_table_591_3_sva <= 1'b0;
      sigmoid_table_591_8_sva <= 1'b0;
      sigmoid_table_590_1_sva <= 1'b0;
      sigmoid_table_590_8_sva <= 1'b0;
      sigmoid_table_589_0_sva <= 1'b0;
      sigmoid_table_589_8_sva <= 1'b0;
      sigmoid_table_588_8_sva <= 1'b0;
      sigmoid_table_587_2_sva <= 1'b0;
      sigmoid_table_587_8_sva <= 1'b0;
      sigmoid_table_586_8_sva <= 1'b0;
      sigmoid_table_585_0_sva <= 1'b0;
      sigmoid_table_585_8_sva <= 1'b0;
      sigmoid_table_584_8_sva <= 1'b0;
      sigmoid_table_583_8_sva <= 1'b0;
      sigmoid_table_582_0_sva <= 1'b0;
      sigmoid_table_581_2_sva <= 1'b0;
      sigmoid_table_580_3_sva <= 1'b0;
      sigmoid_table_579_4_sva <= 1'b0;
      sigmoid_table_578_4_sva <= 1'b0;
      sigmoid_table_577_0_sva <= 1'b0;
      sigmoid_table_577_5_sva <= 1'b0;
      sigmoid_table_576_2_sva <= 1'b0;
      sigmoid_table_576_5_sva <= 1'b0;
      sigmoid_table_575_5_sva <= 1'b0;
      sigmoid_table_574_1_sva <= 1'b0;
      sigmoid_table_574_5_sva <= 1'b0;
      sigmoid_table_573_0_sva <= 1'b0;
      sigmoid_table_573_5_sva <= 1'b0;
      sigmoid_table_572_0_sva <= 1'b0;
      sigmoid_table_572_6_sva <= 1'b0;
      sigmoid_table_571_2_sva <= 1'b0;
      sigmoid_table_571_6_sva <= 1'b0;
      sigmoid_table_570_3_sva <= 1'b0;
      sigmoid_table_570_6_sva <= 1'b0;
      sigmoid_table_569_1_sva <= 1'b0;
      sigmoid_table_569_6_sva <= 1'b0;
      sigmoid_table_568_6_sva <= 1'b0;
      sigmoid_table_567_0_sva <= 1'b0;
      sigmoid_table_567_6_sva <= 1'b0;
      sigmoid_table_566_2_sva <= 1'b0;
      sigmoid_table_566_6_sva <= 1'b0;
      sigmoid_table_565_6_sva <= 1'b0;
      sigmoid_table_564_6_sva <= 1'b0;
      sigmoid_table_563_6_sva <= 1'b0;
      sigmoid_table_562_1_sva <= 1'b0;
      sigmoid_table_561_3_sva <= 1'b0;
      sigmoid_table_560_0_sva <= 1'b0;
      sigmoid_table_560_4_sva <= 1'b0;
      sigmoid_table_559_0_sva <= 1'b0;
      sigmoid_table_559_4_sva <= 1'b0;
      sigmoid_table_558_4_sva <= 1'b0;
      sigmoid_table_557_2_sva <= 1'b0;
      sigmoid_table_553_1_sva <= 1'b0;
      sigmoid_table_552_3_sva <= 1'b0;
      sigmoid_table_551_0_sva <= 1'b0;
      sigmoid_table_550_0_sva <= 1'b0;
      sigmoid_table_548_2_sva <= 1'b0;
      sigmoid_table_544_2_sva <= 1'b0;
      sigmoid_table_543_3_sva <= 1'b0;
      sigmoid_table_542_4_sva <= 1'b0;
      sigmoid_table_541_4_sva <= 1'b0;
      sigmoid_table_540_1_sva <= 1'b0;
      sigmoid_table_540_5_sva <= 1'b0;
      sigmoid_table_539_5_sva <= 1'b0;
      sigmoid_table_538_1_sva <= 1'b0;
      sigmoid_table_538_5_sva <= 1'b0;
      sigmoid_table_537_5_sva <= 1'b0;
      sigmoid_table_536_1_sva <= 1'b0;
      sigmoid_table_535_0_sva <= 1'b0;
      sigmoid_table_535_3_sva <= 1'b0;
      sigmoid_table_534_0_sva <= 1'b0;
      sigmoid_table_533_0_sva <= 1'b0;
      sigmoid_table_532_0_sva <= 1'b0;
      sigmoid_table_531_0_sva <= 1'b0;
      sigmoid_table_530_0_sva <= 1'b0;
      sigmoid_table_529_0_sva <= 1'b0;
      sigmoid_table_528_0_sva <= 1'b0;
      sigmoid_table_527_0_sva <= 1'b0;
      sigmoid_table_527_3_sva <= 1'b0;
      sigmoid_table_526_0_sva <= 1'b0;
      sigmoid_table_526_4_sva <= 1'b0;
      sigmoid_table_525_0_sva <= 1'b0;
      sigmoid_table_525_4_sva <= 1'b0;
      sigmoid_table_524_0_sva <= 1'b0;
      sigmoid_table_523_0_sva <= 1'b0;
      sigmoid_table_522_0_sva <= 1'b0;
      sigmoid_table_521_0_sva <= 1'b0;
      sigmoid_table_520_0_sva <= 1'b0;
      sigmoid_table_519_0_sva <= 1'b0;
      sigmoid_table_519_3_sva <= 1'b0;
      sigmoid_table_518_0_sva <= 1'b0;
      sigmoid_table_517_0_sva <= 1'b0;
      sigmoid_table_516_0_sva <= 1'b0;
      sigmoid_table_515_2_sva <= 1'b0;
      sigmoid_table_511_2_sva <= 1'b0;
      sigmoid_table_510_3_sva <= 1'b0;
      sigmoid_table_509_4_sva <= 1'b0;
      sigmoid_table_508_4_sva <= 1'b0;
      sigmoid_table_507_2_sva <= 1'b0;
      sigmoid_table_507_5_sva <= 1'b0;
      sigmoid_table_506_5_sva <= 1'b0;
      sigmoid_table_505_5_sva <= 1'b0;
      sigmoid_table_504_5_sva <= 1'b0;
      sigmoid_table_503_2_sva <= 1'b0;
      sigmoid_table_503_6_sva <= 1'b0;
      sigmoid_table_502_3_sva <= 1'b0;
      sigmoid_table_502_6_sva <= 1'b0;
      sigmoid_table_501_6_sva <= 1'b0;
      sigmoid_table_500_6_sva <= 1'b0;
      sigmoid_table_499_2_sva <= 1'b0;
      sigmoid_table_499_6_sva <= 1'b0;
      sigmoid_table_498_6_sva <= 1'b0;
      sigmoid_table_497_6_sva <= 1'b0;
      sigmoid_table_496_6_sva <= 1'b0;
      sigmoid_table_495_2_sva <= 1'b0;
      sigmoid_table_495_7_sva <= 1'b0;
      sigmoid_table_494_3_sva <= 1'b0;
      sigmoid_table_494_7_sva <= 1'b0;
      sigmoid_table_493_4_sva <= 1'b0;
      sigmoid_table_493_7_sva <= 1'b0;
      sigmoid_table_492_4_sva <= 1'b0;
      sigmoid_table_492_7_sva <= 1'b0;
      sigmoid_table_491_2_sva <= 1'b0;
      sigmoid_table_491_7_sva <= 1'b0;
      sigmoid_table_490_7_sva <= 1'b0;
      sigmoid_table_489_7_sva <= 1'b0;
      sigmoid_table_488_7_sva <= 1'b0;
      sigmoid_table_487_2_sva <= 1'b0;
      sigmoid_table_487_7_sva <= 1'b0;
      sigmoid_table_486_3_sva <= 1'b0;
      sigmoid_table_486_7_sva <= 1'b0;
      sigmoid_table_485_7_sva <= 1'b0;
      sigmoid_table_484_7_sva <= 1'b0;
      sigmoid_table_483_2_sva <= 1'b0;
      sigmoid_table_483_7_sva <= 1'b0;
      sigmoid_table_482_7_sva <= 1'b0;
      sigmoid_table_481_1_sva <= 1'b0;
      sigmoid_table_481_7_sva <= 1'b0;
      sigmoid_table_480_7_sva <= 1'b0;
      sigmoid_table_479_1_sva <= 1'b0;
      sigmoid_table_478_0_sva <= 1'b0;
      sigmoid_table_478_3_sva <= 1'b0;
      sigmoid_table_477_0_sva <= 1'b0;
      sigmoid_table_477_4_sva <= 1'b0;
      sigmoid_table_476_0_sva <= 1'b0;
      sigmoid_table_476_4_sva <= 1'b0;
      sigmoid_table_475_0_sva <= 1'b0;
      sigmoid_table_475_5_sva <= 1'b0;
      sigmoid_table_474_2_sva <= 1'b0;
      sigmoid_table_474_5_sva <= 1'b0;
      sigmoid_table_473_5_sva <= 1'b0;
      sigmoid_table_472_5_sva <= 1'b0;
      sigmoid_table_471_5_sva <= 1'b0;
      sigmoid_table_470_2_sva <= 1'b0;
      sigmoid_table_469_3_sva <= 1'b0;
      sigmoid_table_468_1_sva <= 1'b0;
      sigmoid_table_467_0_sva <= 1'b0;
      sigmoid_table_466_0_sva <= 1'b0;
      sigmoid_table_465_2_sva <= 1'b0;
      sigmoid_table_461_1_sva <= 1'b0;
      sigmoid_table_460_3_sva <= 1'b0;
      sigmoid_table_459_0_sva <= 1'b0;
      sigmoid_table_459_4_sva <= 1'b0;
      sigmoid_table_458_0_sva <= 1'b0;
      sigmoid_table_458_4_sva <= 1'b0;
      sigmoid_table_457_4_sva <= 1'b0;
      sigmoid_table_456_2_sva <= 1'b0;
      sigmoid_table_454_1_sva <= 1'b0;
      sigmoid_table_453_0_sva <= 1'b0;
      sigmoid_table_451_2_sva <= 1'b0;
      sigmoid_table_450_3_sva <= 1'b0;
      sigmoid_table_449_1_sva <= 1'b0;
      sigmoid_table_448_0_sva <= 1'b0;
      sigmoid_table_446_2_sva <= 1'b0;
      sigmoid_table_444_1_sva <= 1'b0;
      sigmoid_table_443_0_sva <= 1'b0;
      sigmoid_table_441_2_sva <= 1'b0;
      sigmoid_table_440_3_sva <= 1'b0;
      sigmoid_table_439_3_sva <= 1'b0;
      sigmoid_table_438_4_sva <= 1'b0;
      sigmoid_table_437_4_sva <= 1'b0;
      sigmoid_table_436_0_sva <= 1'b0;
      sigmoid_table_436_5_sva <= 1'b0;
      sigmoid_table_435_2_sva <= 1'b0;
      sigmoid_table_435_5_sva <= 1'b0;
      sigmoid_table_434_5_sva <= 1'b0;
      sigmoid_table_433_1_sva <= 1'b0;
      sigmoid_table_433_5_sva <= 1'b0;
      sigmoid_table_432_5_sva <= 1'b0;
      sigmoid_table_431_5_sva <= 1'b0;
      sigmoid_table_430_1_sva <= 1'b0;
      sigmoid_table_430_6_sva <= 1'b0;
      sigmoid_table_429_0_sva <= 1'b0;
      sigmoid_table_429_3_sva <= 1'b0;
      sigmoid_table_429_6_sva <= 1'b0;
      sigmoid_table_428_3_sva <= 1'b0;
      sigmoid_table_428_6_sva <= 1'b0;
      sigmoid_table_427_1_sva <= 1'b0;
      sigmoid_table_427_6_sva <= 1'b0;
      sigmoid_table_426_0_sva <= 1'b0;
      sigmoid_table_426_6_sva <= 1'b0;
      sigmoid_table_425_6_sva <= 1'b0;
      sigmoid_table_424_1_sva <= 1'b0;
      sigmoid_table_424_6_sva <= 1'b0;
      sigmoid_table_423_2_sva <= 1'b0;
      sigmoid_table_423_6_sva <= 1'b0;
      sigmoid_table_422_6_sva <= 1'b0;
      sigmoid_table_421_0_sva <= 1'b0;
      sigmoid_table_421_6_sva <= 1'b0;
      sigmoid_table_420_6_sva <= 1'b0;
      sigmoid_table_419_6_sva <= 1'b0;
      sigmoid_table_418_0_sva <= 1'b0;
      sigmoid_table_417_2_sva <= 1'b0;
      sigmoid_table_416_3_sva <= 1'b0;
      sigmoid_table_415_3_sva <= 1'b0;
      sigmoid_table_414_1_sva <= 1'b0;
      sigmoid_table_414_4_sva <= 1'b0;
      sigmoid_table_413_0_sva <= 1'b0;
      sigmoid_table_413_4_sva <= 1'b0;
      sigmoid_table_412_4_sva <= 1'b0;
      sigmoid_table_411_0_sva <= 1'b0;
      sigmoid_table_410_2_sva <= 1'b0;
      sigmoid_table_407_1_sva <= 1'b0;
      sigmoid_table_404_0_sva <= 1'b0;
      sigmoid_table_403_2_sva <= 1'b0;
      sigmoid_table_402_0_sva <= 1'b0;
      sigmoid_table_402_3_sva <= 1'b0;
      sigmoid_table_401_3_sva <= 1'b0;
      sigmoid_table_400_0_sva <= 1'b0;
      sigmoid_table_398_0_sva <= 1'b0;
      sigmoid_table_396_0_sva <= 1'b0;
      sigmoid_table_395_2_sva <= 1'b0;
      sigmoid_table_394_0_sva <= 1'b0;
      sigmoid_table_391_1_sva <= 1'b0;
      sigmoid_table_387_0_sva <= 1'b0;
      sigmoid_table_386_2_sva <= 1'b0;
      sigmoid_table_385_0_sva <= 1'b0;
      sigmoid_table_385_3_sva <= 1'b0;
      sigmoid_table_384_3_sva <= 1'b0;
      sigmoid_table_383_3_sva <= 1'b0;
      sigmoid_table_382_1_sva <= 1'b0;
      sigmoid_table_382_4_sva <= 1'b0;
      sigmoid_table_381_4_sva <= 1'b0;
      sigmoid_table_380_0_sva <= 1'b0;
      sigmoid_table_380_4_sva <= 1'b0;
      sigmoid_table_379_4_sva <= 1'b0;
      sigmoid_table_378_4_sva <= 1'b0;
      sigmoid_table_377_1_sva <= 1'b0;
      sigmoid_table_377_5_sva <= 1'b0;
      sigmoid_table_376_2_sva <= 1'b0;
      sigmoid_table_376_5_sva <= 1'b0;
      sigmoid_table_375_0_sva <= 1'b0;
      sigmoid_table_375_5_sva <= 1'b0;
      sigmoid_table_374_5_sva <= 1'b0;
      sigmoid_table_373_5_sva <= 1'b0;
      sigmoid_table_372_0_sva <= 1'b0;
      sigmoid_table_372_5_sva <= 1'b0;
      sigmoid_table_371_5_sva <= 1'b0;
      sigmoid_table_370_5_sva <= 1'b0;
      sigmoid_table_369_0_sva <= 1'b0;
      sigmoid_table_369_5_sva <= 1'b0;
      sigmoid_table_368_5_sva <= 1'b0;
      sigmoid_table_367_5_sva <= 1'b0;
      sigmoid_table_366_1_sva <= 1'b0;
      sigmoid_table_365_2_sva <= 1'b0;
      sigmoid_table_364_2_sva <= 1'b0;
      sigmoid_table_363_3_sva <= 1'b0;
      sigmoid_table_362_3_sva <= 1'b0;
      sigmoid_table_361_3_sva <= 1'b0;
      sigmoid_table_360_0_sva <= 1'b0;
      sigmoid_table_357_0_sva <= 1'b0;
      sigmoid_table_354_0_sva <= 1'b0;
      sigmoid_table_353_1_sva <= 1'b0;
      sigmoid_table_352_2_sva <= 1'b0;
      sigmoid_table_351_2_sva <= 1'b0;
      sigmoid_table_350_0_sva <= 1'b0;
      sigmoid_table_346_0_sva <= 1'b0;
      sigmoid_table_345_1_sva <= 1'b0;
      sigmoid_table_342_0_sva <= 1'b0;
      sigmoid_table_338_0_sva <= 1'b0;
      sigmoid_table_337_1_sva <= 1'b0;
      sigmoid_table_336_2_sva <= 1'b0;
      sigmoid_table_335_2_sva <= 1'b0;
      sigmoid_table_334_0_sva <= 1'b0;
      sigmoid_table_334_3_sva <= 1'b0;
      sigmoid_table_333_3_sva <= 1'b0;
      sigmoid_table_332_3_sva <= 1'b0;
      sigmoid_table_331_3_sva <= 1'b0;
      sigmoid_table_330_3_sva <= 1'b0;
      sigmoid_table_329_0_sva <= 1'b0;
      sigmoid_table_329_4_sva <= 1'b0;
      sigmoid_table_328_1_sva <= 1'b0;
      sigmoid_table_328_4_sva <= 1'b0;
      sigmoid_table_327_4_sva <= 1'b0;
      sigmoid_table_326_4_sva <= 1'b0;
      sigmoid_table_325_4_sva <= 1'b0;
      sigmoid_table_324_0_sva <= 1'b0;
      sigmoid_table_324_4_sva <= 1'b0;
      sigmoid_table_323_4_sva <= 1'b0;
      sigmoid_table_322_4_sva <= 1'b0;
      sigmoid_table_321_4_sva <= 1'b0;
      sigmoid_table_320_4_sva <= 1'b0;
      sigmoid_table_319_0_sva <= 1'b0;
      sigmoid_table_318_0_sva <= 1'b0;
      sigmoid_table_317_1_sva <= 1'b0;
      sigmoid_table_316_2_sva <= 1'b0;
      sigmoid_table_315_2_sva <= 1'b0;
      sigmoid_table_314_2_sva <= 1'b0;
      sigmoid_table_313_0_sva <= 1'b0;
      sigmoid_table_312_0_sva <= 1'b0;
      sigmoid_table_307_0_sva <= 1'b0;
      sigmoid_table_306_0_sva <= 1'b0;
      sigmoid_table_305_1_sva <= 1'b0;
      sigmoid_table_304_1_sva <= 1'b0;
      sigmoid_table_300_0_sva <= 1'b0;
      sigmoid_table_299_0_sva <= 1'b0;
      sigmoid_table_292_0_sva <= 1'b0;
      sigmoid_table_291_0_sva <= 1'b0;
      sigmoid_table_290_1_sva <= 1'b0;
      sigmoid_table_289_1_sva <= 1'b0;
      sigmoid_table_288_1_sva <= 1'b0;
      sigmoid_table_287_2_sva <= 1'b0;
      sigmoid_table_286_2_sva <= 1'b0;
      sigmoid_table_285_2_sva <= 1'b0;
      sigmoid_table_284_2_sva <= 1'b0;
      sigmoid_table_283_0_sva <= 1'b0;
      sigmoid_table_283_3_sva <= 1'b0;
      sigmoid_table_282_0_sva <= 1'b0;
      sigmoid_table_282_3_sva <= 1'b0;
      sigmoid_table_281_3_sva <= 1'b0;
      sigmoid_table_280_3_sva <= 1'b0;
      sigmoid_table_279_3_sva <= 1'b0;
      sigmoid_table_278_3_sva <= 1'b0;
      sigmoid_table_277_3_sva <= 1'b0;
      sigmoid_table_276_3_sva <= 1'b0;
      sigmoid_table_275_3_sva <= 1'b0;
      sigmoid_table_274_3_sva <= 1'b0;
      sigmoid_table_273_0_sva <= 1'b0;
      sigmoid_table_272_0_sva <= 1'b0;
      sigmoid_table_271_0_sva <= 1'b0;
      sigmoid_table_270_1_sva <= 1'b0;
      sigmoid_table_269_1_sva <= 1'b0;
      sigmoid_table_268_1_sva <= 1'b0;
      sigmoid_table_261_0_sva <= 1'b0;
      sigmoid_table_260_0_sva <= 1'b0;
      sigmoid_table_259_0_sva <= 1'b0;
      sigmoid_table_246_0_sva <= 1'b0;
      sigmoid_table_245_0_sva <= 1'b0;
      sigmoid_table_244_0_sva <= 1'b0;
      sigmoid_table_243_0_sva <= 1'b0;
      sigmoid_table_242_1_sva <= 1'b0;
      sigmoid_table_241_1_sva <= 1'b0;
      sigmoid_table_240_1_sva <= 1'b0;
      sigmoid_table_239_1_sva <= 1'b0;
      sigmoid_table_238_2_sva <= 1'b0;
      sigmoid_table_237_2_sva <= 1'b0;
      sigmoid_table_236_2_sva <= 1'b0;
      sigmoid_table_235_2_sva <= 1'b0;
      sigmoid_table_234_2_sva <= 1'b0;
      sigmoid_table_233_2_sva <= 1'b0;
      sigmoid_table_232_2_sva <= 1'b0;
      sigmoid_table_231_2_sva <= 1'b0;
      sigmoid_table_230_2_sva <= 1'b0;
      sigmoid_table_229_2_sva <= 1'b0;
      sigmoid_table_228_0_sva <= 1'b0;
      sigmoid_table_227_0_sva <= 1'b0;
      sigmoid_table_226_0_sva <= 1'b0;
      sigmoid_table_225_0_sva <= 1'b0;
      sigmoid_table_224_0_sva <= 1'b0;
      sigmoid_table_223_0_sva <= 1'b0;
      sigmoid_table_201_0_sva <= 1'b0;
      sigmoid_table_200_0_sva <= 1'b0;
      sigmoid_table_199_0_sva <= 1'b0;
      sigmoid_table_198_0_sva <= 1'b0;
      sigmoid_table_197_0_sva <= 1'b0;
      sigmoid_table_196_0_sva <= 1'b0;
      sigmoid_table_195_0_sva <= 1'b0;
      sigmoid_table_194_0_sva <= 1'b0;
      sigmoid_table_193_1_sva <= 1'b0;
      sigmoid_table_192_1_sva <= 1'b0;
      sigmoid_table_191_1_sva <= 1'b0;
      sigmoid_table_190_1_sva <= 1'b0;
      sigmoid_table_189_1_sva <= 1'b0;
      sigmoid_table_188_1_sva <= 1'b0;
      sigmoid_table_187_1_sva <= 1'b0;
      sigmoid_table_186_1_sva <= 1'b0;
      sigmoid_table_185_1_sva <= 1'b0;
      sigmoid_table_184_1_sva <= 1'b0;
      sigmoid_table_157_0_sva <= 1'b0;
      sigmoid_table_156_0_sva <= 1'b0;
      sigmoid_table_155_0_sva <= 1'b0;
      sigmoid_table_154_0_sva <= 1'b0;
      sigmoid_table_153_0_sva <= 1'b0;
      sigmoid_table_152_0_sva <= 1'b0;
      sigmoid_table_151_0_sva <= 1'b0;
      sigmoid_table_150_0_sva <= 1'b0;
      sigmoid_table_149_0_sva <= 1'b0;
      sigmoid_table_148_0_sva <= 1'b0;
      sigmoid_table_147_0_sva <= 1'b0;
      sigmoid_table_146_0_sva <= 1'b0;
      sigmoid_table_145_0_sva <= 1'b0;
      sigmoid_table_144_0_sva <= 1'b0;
      sigmoid_table_143_0_sva <= 1'b0;
      sigmoid_table_142_0_sva <= 1'b0;
      sigmoid_table_141_0_sva <= 1'b0;
      sigmoid_table_140_0_sva <= 1'b0;
      sigmoid_table_139_0_sva <= 1'b0;
      sigmoid_table_910_0_sva <= 1'b0;
      sigmoid_table_909_0_sva <= 1'b0;
      sigmoid_table_908_0_sva <= 1'b0;
      sigmoid_table_907_0_sva <= 1'b0;
      sigmoid_table_906_0_sva <= 1'b0;
      sigmoid_table_905_0_sva <= 1'b0;
      sigmoid_table_904_0_sva <= 1'b0;
      sigmoid_table_903_0_sva <= 1'b0;
      sigmoid_table_902_0_sva <= 1'b0;
      sigmoid_table_901_0_sva <= 1'b0;
      sigmoid_table_900_0_sva <= 1'b0;
      sigmoid_table_899_0_sva <= 1'b0;
      sigmoid_table_898_0_sva <= 1'b0;
      sigmoid_table_897_0_sva <= 1'b0;
      sigmoid_table_896_0_sva <= 1'b0;
      sigmoid_table_895_0_sva <= 1'b0;
      sigmoid_table_894_0_sva <= 1'b0;
      sigmoid_table_893_0_sva <= 1'b0;
      sigmoid_table_892_0_sva <= 1'b0;
      sigmoid_table_891_0_sva <= 1'b0;
      sigmoid_table_890_0_sva <= 1'b0;
      sigmoid_table_889_0_sva <= 1'b0;
      sigmoid_table_888_0_sva <= 1'b0;
      sigmoid_table_887_0_sva <= 1'b0;
      sigmoid_table_886_0_sva <= 1'b0;
      sigmoid_table_885_0_sva <= 1'b0;
      sigmoid_table_852_1_sva <= 1'b0;
      sigmoid_table_851_1_sva <= 1'b0;
      sigmoid_table_850_1_sva <= 1'b0;
      sigmoid_table_849_1_sva <= 1'b0;
      sigmoid_table_848_1_sva <= 1'b0;
      sigmoid_table_847_1_sva <= 1'b0;
      sigmoid_table_846_1_sva <= 1'b0;
      sigmoid_table_845_1_sva <= 1'b0;
      sigmoid_table_844_1_sva <= 1'b0;
      sigmoid_table_843_1_sva <= 1'b0;
      sigmoid_table_842_1_sva <= 1'b0;
      sigmoid_table_841_1_sva <= 1'b0;
      sigmoid_table_840_0_sva <= 1'b0;
      sigmoid_table_839_0_sva <= 1'b0;
      sigmoid_table_838_0_sva <= 1'b0;
      sigmoid_table_837_0_sva <= 1'b0;
      sigmoid_table_836_0_sva <= 1'b0;
      sigmoid_table_835_0_sva <= 1'b0;
      sigmoid_table_834_0_sva <= 1'b0;
      sigmoid_table_833_0_sva <= 1'b0;
      sigmoid_table_832_0_sva <= 1'b0;
      sigmoid_table_831_0_sva <= 1'b0;
      sigmoid_table_807_0_sva <= 1'b0;
      sigmoid_table_807_2_sva <= 1'b0;
      sigmoid_table_806_0_sva <= 1'b0;
      sigmoid_table_806_2_sva <= 1'b0;
      sigmoid_table_805_0_sva <= 1'b0;
      sigmoid_table_805_2_sva <= 1'b0;
      sigmoid_table_804_0_sva <= 1'b0;
      sigmoid_table_804_2_sva <= 1'b0;
      sigmoid_table_803_0_sva <= 1'b0;
      sigmoid_table_803_2_sva <= 1'b0;
      sigmoid_table_802_0_sva <= 1'b0;
      sigmoid_table_802_2_sva <= 1'b0;
      sigmoid_table_801_2_sva <= 1'b0;
      sigmoid_table_800_2_sva <= 1'b0;
      sigmoid_table_799_2_sva <= 1'b0;
      sigmoid_table_798_2_sva <= 1'b0;
      sigmoid_table_797_2_sva <= 1'b0;
      sigmoid_table_796_2_sva <= 1'b0;
      sigmoid_table_790_1_sva <= 1'b0;
      sigmoid_table_789_1_sva <= 1'b0;
      sigmoid_table_788_1_sva <= 1'b0;
      sigmoid_table_787_1_sva <= 1'b0;
      sigmoid_table_786_1_sva <= 1'b0;
      sigmoid_table_785_0_sva <= 1'b0;
      sigmoid_table_784_0_sva <= 1'b0;
      sigmoid_table_783_0_sva <= 1'b0;
      sigmoid_table_782_0_sva <= 1'b0;
      sigmoid_table_769_0_sva <= 1'b0;
      sigmoid_table_768_0_sva <= 1'b0;
      sigmoid_table_767_0_sva <= 1'b0;
      sigmoid_table_766_0_sva <= 1'b0;
      sigmoid_table_762_3_sva <= 1'b0;
      sigmoid_table_761_3_sva <= 1'b0;
      sigmoid_table_760_3_sva <= 1'b0;
      sigmoid_table_759_1_sva <= 1'b0;
      sigmoid_table_759_3_sva <= 1'b0;
      sigmoid_table_758_1_sva <= 1'b0;
      sigmoid_table_758_3_sva <= 1'b0;
      sigmoid_table_757_1_sva <= 1'b0;
      sigmoid_table_757_3_sva <= 1'b0;
      sigmoid_table_756_0_sva <= 1'b0;
      sigmoid_table_756_3_sva <= 1'b0;
      sigmoid_table_755_0_sva <= 1'b0;
      sigmoid_table_755_3_sva <= 1'b0;
      sigmoid_table_754_0_sva <= 1'b0;
      sigmoid_table_754_3_sva <= 1'b0;
      sigmoid_table_753_3_sva <= 1'b0;
      sigmoid_table_752_3_sva <= 1'b0;
      sigmoid_table_751_3_sva <= 1'b0;
      sigmoid_table_745_0_sva <= 1'b0;
      sigmoid_table_745_2_sva <= 1'b0;
      sigmoid_table_744_0_sva <= 1'b0;
      sigmoid_table_744_2_sva <= 1'b0;
      sigmoid_table_743_0_sva <= 1'b0;
      sigmoid_table_743_2_sva <= 1'b0;
      sigmoid_table_742_2_sva <= 1'b0;
      sigmoid_table_741_2_sva <= 1'b0;
      sigmoid_table_738_1_sva <= 1'b0;
      sigmoid_table_737_1_sva <= 1'b0;
      sigmoid_table_736_0_sva <= 1'b0;
      sigmoid_table_735_0_sva <= 1'b0;
      sigmoid_table_734_0_sva <= 1'b0;
      sigmoid_table_727_0_sva <= 1'b0;
      sigmoid_table_726_0_sva <= 1'b0;
      sigmoid_table_722_1_sva <= 1'b0;
      sigmoid_table_721_1_sva <= 1'b0;
      sigmoid_table_720_0_sva <= 1'b0;
      sigmoid_table_719_0_sva <= 1'b0;
      sigmoid_table_716_4_sva <= 1'b0;
      sigmoid_table_715_4_sva <= 1'b0;
      sigmoid_table_714_4_sva <= 1'b0;
      sigmoid_table_713_0_sva <= 1'b0;
      sigmoid_table_713_2_sva <= 1'b0;
      sigmoid_table_713_4_sva <= 1'b0;
      sigmoid_table_712_2_sva <= 1'b0;
      sigmoid_table_712_4_sva <= 1'b0;
      sigmoid_table_711_2_sva <= 1'b0;
      sigmoid_table_711_4_sva <= 1'b0;
      sigmoid_table_710_4_sva <= 1'b0;
      sigmoid_table_709_1_sva <= 1'b0;
      sigmoid_table_709_4_sva <= 1'b0;
      sigmoid_table_708_1_sva <= 1'b0;
      sigmoid_table_708_4_sva <= 1'b0;
      sigmoid_table_707_0_sva <= 1'b0;
      sigmoid_table_707_4_sva <= 1'b0;
      sigmoid_table_706_4_sva <= 1'b0;
      sigmoid_table_705_4_sva <= 1'b0;
      sigmoid_table_702_0_sva <= 1'b0;
      sigmoid_table_701_0_sva <= 1'b0;
      sigmoid_table_699_3_sva <= 1'b0;
      sigmoid_table_698_1_sva <= 1'b0;
      sigmoid_table_698_3_sva <= 1'b0;
      sigmoid_table_697_1_sva <= 1'b0;
      sigmoid_table_697_3_sva <= 1'b0;
      sigmoid_table_696_0_sva <= 1'b0;
      sigmoid_table_696_3_sva <= 1'b0;
      sigmoid_table_695_3_sva <= 1'b0;
      sigmoid_table_692_0_sva <= 1'b0;
      sigmoid_table_692_2_sva <= 1'b0;
      sigmoid_table_691_0_sva <= 1'b0;
      sigmoid_table_691_2_sva <= 1'b0;
      sigmoid_table_690_2_sva <= 1'b0;
      sigmoid_table_688_1_sva <= 1'b0;
      sigmoid_table_687_0_sva <= 1'b0;
      sigmoid_table_683_0_sva <= 1'b0;
      sigmoid_table_680_1_sva <= 1'b0;
      sigmoid_table_679_0_sva <= 1'b0;
      sigmoid_table_675_0_sva <= 1'b0;
      sigmoid_table_675_2_sva <= 1'b0;
      sigmoid_table_674_2_sva <= 1'b0;
      sigmoid_table_672_1_sva <= 1'b0;
      sigmoid_table_671_0_sva <= 1'b0;
      sigmoid_table_669_5_sva <= 1'b0;
      sigmoid_table_668_0_sva <= 1'b0;
      sigmoid_table_668_5_sva <= 1'b0;
      sigmoid_table_667_5_sva <= 1'b0;
      sigmoid_table_666_3_sva <= 1'b0;
      sigmoid_table_666_5_sva <= 1'b0;
      sigmoid_table_665_1_sva <= 1'b0;
      sigmoid_table_665_3_sva <= 1'b0;
      sigmoid_table_665_5_sva <= 1'b0;
      sigmoid_table_664_3_sva <= 1'b0;
      sigmoid_table_664_5_sva <= 1'b0;
      sigmoid_table_663_5_sva <= 1'b0;
      sigmoid_table_662_5_sva <= 1'b0;
      sigmoid_table_661_0_sva <= 1'b0;
      sigmoid_table_661_2_sva <= 1'b0;
      sigmoid_table_661_5_sva <= 1'b0;
      sigmoid_table_660_5_sva <= 1'b0;
      sigmoid_table_659_1_sva <= 1'b0;
      sigmoid_table_659_5_sva <= 1'b0;
      sigmoid_table_658_0_sva <= 1'b0;
      sigmoid_table_658_5_sva <= 1'b0;
      sigmoid_table_653_1_sva <= 1'b0;
      sigmoid_table_651_4_sva <= 1'b0;
      sigmoid_table_650_0_sva <= 1'b0;
      sigmoid_table_650_2_sva <= 1'b0;
      sigmoid_table_650_4_sva <= 1'b0;
      sigmoid_table_649_2_sva <= 1'b0;
      sigmoid_table_649_4_sva <= 1'b0;
      sigmoid_table_648_1_sva <= 1'b0;
      sigmoid_table_648_4_sva <= 1'b0;
      sigmoid_table_647_0_sva <= 1'b0;
      sigmoid_table_647_4_sva <= 1'b0;
      sigmoid_table_643_1_sva <= 1'b0;
      sigmoid_table_643_3_sva <= 1'b0;
      sigmoid_table_642_0_sva <= 1'b0;
      sigmoid_table_642_3_sva <= 1'b0;
      sigmoid_table_640_0_sva <= 1'b0;
      sigmoid_table_640_2_sva <= 1'b0;
      sigmoid_table_639_2_sva <= 1'b0;
      sigmoid_table_638_1_sva <= 1'b0;
      sigmoid_table_635_0_sva <= 1'b0;
      sigmoid_table_633_0_sva <= 1'b0;
      sigmoid_table_631_0_sva <= 1'b0;
      sigmoid_table_631_2_sva <= 1'b0;
      sigmoid_table_630_2_sva <= 1'b0;
      sigmoid_table_629_1_sva <= 1'b0;
      sigmoid_table_625_1_sva <= 1'b0;
      sigmoid_table_625_3_sva <= 1'b0;
      sigmoid_table_624_3_sva <= 1'b0;
      sigmoid_table_622_2_sva <= 1'b0;
      sigmoid_table_621_1_sva <= 1'b0;
      sigmoid_table_619_6_sva <= 1'b0;
      sigmoid_table_618_6_sva <= 1'b0;
      sigmoid_table_617_0_sva <= 1'b0;
      sigmoid_table_617_6_sva <= 1'b0;
      sigmoid_table_616_4_sva <= 1'b0;
      sigmoid_table_616_6_sva <= 1'b0;
      sigmoid_table_615_0_sva <= 1'b0;
      sigmoid_table_615_2_sva <= 1'b0;
      sigmoid_table_615_4_sva <= 1'b0;
      sigmoid_table_615_6_sva <= 1'b0;
      sigmoid_table_614_4_sva <= 1'b0;
      sigmoid_table_614_6_sva <= 1'b0;
      sigmoid_table_613_4_sva <= 1'b0;
      sigmoid_table_613_6_sva <= 1'b0;
      sigmoid_table_612_6_sva <= 1'b0;
      sigmoid_table_611_6_sva <= 1'b0;
      sigmoid_table_610_0_sva <= 1'b0;
      sigmoid_table_610_3_sva <= 1'b0;
      sigmoid_table_610_6_sva <= 1'b0;
      sigmoid_table_609_6_sva <= 1'b0;
      sigmoid_table_608_0_sva <= 1'b0;
      sigmoid_table_608_2_sva <= 1'b0;
      sigmoid_table_608_6_sva <= 1'b0;
      sigmoid_table_607_1_sva <= 1'b0;
      sigmoid_table_607_6_sva <= 1'b0;
      sigmoid_table_606_6_sva <= 1'b0;
      sigmoid_table_605_0_sva <= 1'b0;
      sigmoid_table_600_0_sva <= 1'b0;
      sigmoid_table_599_5_sva <= 1'b0;
      sigmoid_table_598_5_sva <= 1'b0;
      sigmoid_table_597_0_sva <= 1'b0;
      sigmoid_table_597_3_sva <= 1'b0;
      sigmoid_table_597_5_sva <= 1'b0;
      sigmoid_table_596_5_sva <= 1'b0;
      sigmoid_table_595_2_sva <= 1'b0;
      sigmoid_table_595_5_sva <= 1'b0;
      sigmoid_table_594_0_sva <= 1'b0;
      sigmoid_table_594_5_sva <= 1'b0;
      sigmoid_table_591_0_sva <= 1'b0;
      sigmoid_table_590_4_sva <= 1'b0;
      sigmoid_table_589_4_sva <= 1'b0;
      sigmoid_table_588_4_sva <= 1'b0;
      sigmoid_table_587_0_sva <= 1'b0;
      sigmoid_table_586_1_sva <= 1'b0;
      sigmoid_table_586_3_sva <= 1'b0;
      sigmoid_table_584_0_sva <= 1'b0;
      sigmoid_table_584_2_sva <= 1'b0;
      sigmoid_table_583_1_sva <= 1'b0;
      sigmoid_table_582_9_sva <= 1'b0;
      sigmoid_table_581_9_sva <= 1'b0;
      sigmoid_table_580_0_sva <= 1'b0;
      sigmoid_table_580_9_sva <= 1'b0;
      sigmoid_table_579_0_sva <= 1'b0;
      sigmoid_table_579_2_sva <= 1'b0;
      sigmoid_table_579_9_sva <= 1'b0;
      sigmoid_table_578_1_sva <= 1'b0;
      sigmoid_table_578_9_sva <= 1'b0;
      sigmoid_table_577_9_sva <= 1'b0;
      sigmoid_table_576_9_sva <= 1'b0;
      sigmoid_table_575_0_sva <= 1'b0;
      sigmoid_table_575_3_sva <= 1'b0;
      sigmoid_table_575_9_sva <= 1'b0;
      sigmoid_table_574_9_sva <= 1'b0;
      sigmoid_table_573_9_sva <= 1'b0;
      sigmoid_table_572_9_sva <= 1'b0;
      sigmoid_table_571_9_sva <= 1'b0;
      sigmoid_table_570_0_sva <= 1'b0;
      sigmoid_table_570_9_sva <= 1'b0;
      sigmoid_table_569_4_sva <= 1'b0;
      sigmoid_table_569_9_sva <= 1'b0;
      sigmoid_table_568_1_sva <= 1'b0;
      sigmoid_table_568_4_sva <= 1'b0;
      sigmoid_table_568_9_sva <= 1'b0;
      sigmoid_table_567_9_sva <= 1'b0;
      sigmoid_table_566_9_sva <= 1'b0;
      sigmoid_table_565_3_sva <= 1'b0;
      sigmoid_table_565_9_sva <= 1'b0;
      sigmoid_table_564_0_sva <= 1'b0;
      sigmoid_table_564_2_sva <= 1'b0;
      sigmoid_table_564_9_sva <= 1'b0;
      sigmoid_table_563_0_sva <= 1'b0;
      sigmoid_table_563_9_sva <= 1'b0;
      sigmoid_table_562_7_sva <= 1'b0;
      sigmoid_table_562_9_sva <= 1'b0;
      sigmoid_table_561_1_sva <= 1'b0;
      sigmoid_table_561_7_sva <= 1'b0;
      sigmoid_table_561_9_sva <= 1'b0;
      sigmoid_table_560_7_sva <= 1'b0;
      sigmoid_table_560_9_sva <= 1'b0;
      sigmoid_table_559_7_sva <= 1'b0;
      sigmoid_table_559_9_sva <= 1'b0;
      sigmoid_table_558_7_sva <= 1'b0;
      sigmoid_table_558_9_sva <= 1'b0;
      sigmoid_table_557_5_sva <= 1'b0;
      sigmoid_table_557_7_sva <= 1'b0;
      sigmoid_table_557_9_sva <= 1'b0;
      sigmoid_table_556_0_sva <= 1'b0;
      sigmoid_table_556_3_sva <= 1'b0;
      sigmoid_table_556_5_sva <= 1'b0;
      sigmoid_table_556_7_sva <= 1'b0;
      sigmoid_table_556_9_sva <= 1'b0;
      sigmoid_table_555_0_sva <= 1'b0;
      sigmoid_table_555_2_sva <= 1'b0;
      sigmoid_table_555_5_sva <= 1'b0;
      sigmoid_table_555_7_sva <= 1'b0;
      sigmoid_table_555_9_sva <= 1'b0;
      sigmoid_table_554_1_sva <= 1'b0;
      sigmoid_table_554_5_sva <= 1'b0;
      sigmoid_table_554_7_sva <= 1'b0;
      sigmoid_table_554_9_sva <= 1'b0;
      sigmoid_table_553_7_sva <= 1'b0;
      sigmoid_table_553_9_sva <= 1'b0;
      sigmoid_table_552_1_sva <= 1'b0;
      sigmoid_table_552_7_sva <= 1'b0;
      sigmoid_table_552_9_sva <= 1'b0;
      sigmoid_table_551_4_sva <= 1'b0;
      sigmoid_table_551_7_sva <= 1'b0;
      sigmoid_table_551_9_sva <= 1'b0;
      sigmoid_table_550_4_sva <= 1'b0;
      sigmoid_table_550_7_sva <= 1'b0;
      sigmoid_table_550_9_sva <= 1'b0;
      sigmoid_table_549_4_sva <= 1'b0;
      sigmoid_table_549_7_sva <= 1'b0;
      sigmoid_table_549_9_sva <= 1'b0;
      sigmoid_table_548_7_sva <= 1'b0;
      sigmoid_table_548_9_sva <= 1'b0;
      sigmoid_table_547_3_sva <= 1'b0;
      sigmoid_table_547_7_sva <= 1'b0;
      sigmoid_table_547_9_sva <= 1'b0;
      sigmoid_table_546_2_sva <= 1'b0;
      sigmoid_table_546_7_sva <= 1'b0;
      sigmoid_table_546_9_sva <= 1'b0;
      sigmoid_table_545_0_sva <= 1'b0;
      sigmoid_table_545_7_sva <= 1'b0;
      sigmoid_table_545_9_sva <= 1'b0;
      sigmoid_table_544_0_sva <= 1'b0;
      sigmoid_table_544_9_sva <= 1'b0;
      sigmoid_table_543_0_sva <= 1'b0;
      sigmoid_table_543_9_sva <= 1'b0;
      sigmoid_table_542_0_sva <= 1'b0;
      sigmoid_table_542_2_sva <= 1'b0;
      sigmoid_table_542_9_sva <= 1'b0;
      sigmoid_table_541_1_sva <= 1'b0;
      sigmoid_table_541_9_sva <= 1'b0;
      sigmoid_table_540_9_sva <= 1'b0;
      sigmoid_table_539_1_sva <= 1'b0;
      sigmoid_table_539_3_sva <= 1'b0;
      sigmoid_table_539_9_sva <= 1'b0;
      sigmoid_table_538_9_sva <= 1'b0;
      sigmoid_table_537_1_sva <= 1'b0;
      sigmoid_table_537_9_sva <= 1'b0;
      sigmoid_table_536_6_sva <= 1'b0;
      sigmoid_table_536_9_sva <= 1'b0;
      sigmoid_table_535_6_sva <= 1'b0;
      sigmoid_table_535_9_sva <= 1'b0;
      sigmoid_table_534_4_sva <= 1'b0;
      sigmoid_table_534_6_sva <= 1'b0;
      sigmoid_table_534_9_sva <= 1'b0;
      sigmoid_table_533_4_sva <= 1'b0;
      sigmoid_table_533_6_sva <= 1'b0;
      sigmoid_table_533_9_sva <= 1'b0;
      sigmoid_table_532_6_sva <= 1'b0;
      sigmoid_table_532_9_sva <= 1'b0;
      sigmoid_table_531_3_sva <= 1'b0;
      sigmoid_table_531_6_sva <= 1'b0;
      sigmoid_table_531_9_sva <= 1'b0;
      sigmoid_table_530_6_sva <= 1'b0;
      sigmoid_table_530_9_sva <= 1'b0;
      sigmoid_table_529_6_sva <= 1'b0;
      sigmoid_table_529_9_sva <= 1'b0;
      sigmoid_table_528_9_sva <= 1'b0;
      sigmoid_table_527_9_sva <= 1'b0;
      sigmoid_table_526_9_sva <= 1'b0;
      sigmoid_table_525_9_sva <= 1'b0;
      sigmoid_table_524_5_sva <= 1'b0;
      sigmoid_table_524_9_sva <= 1'b0;
      sigmoid_table_523_3_sva <= 1'b0;
      sigmoid_table_523_5_sva <= 1'b0;
      sigmoid_table_523_9_sva <= 1'b0;
      sigmoid_table_522_5_sva <= 1'b0;
      sigmoid_table_522_9_sva <= 1'b0;
      sigmoid_table_521_5_sva <= 1'b0;
      sigmoid_table_521_9_sva <= 1'b0;
      sigmoid_table_520_9_sva <= 1'b0;
      sigmoid_table_519_9_sva <= 1'b0;
      sigmoid_table_518_4_sva <= 1'b0;
      sigmoid_table_518_9_sva <= 1'b0;
      sigmoid_table_517_4_sva <= 1'b0;
      sigmoid_table_517_9_sva <= 1'b0;
      sigmoid_table_516_9_sva <= 1'b0;
      sigmoid_table_515_9_sva <= 1'b0;
      sigmoid_table_514_3_sva <= 1'b0;
      sigmoid_table_514_9_sva <= 1'b0;
      sigmoid_table_513_2_sva <= 1'b0;
      sigmoid_table_513_9_sva <= 1'b0;
      sigmoid_table_512_9_sva <= 1'b0;
      sigmoid_table_509_2_sva <= 1'b0;
      sigmoid_table_506_3_sva <= 1'b0;
      sigmoid_table_505_2_sva <= 1'b0;
      sigmoid_table_501_2_sva <= 1'b0;
      sigmoid_table_501_4_sva <= 1'b0;
      sigmoid_table_500_4_sva <= 1'b0;
      sigmoid_table_498_3_sva <= 1'b0;
      sigmoid_table_497_2_sva <= 1'b0;
      sigmoid_table_493_2_sva <= 1'b0;
      sigmoid_table_491_5_sva <= 1'b0;
      sigmoid_table_490_3_sva <= 1'b0;
      sigmoid_table_490_5_sva <= 1'b0;
      sigmoid_table_489_2_sva <= 1'b0;
      sigmoid_table_489_5_sva <= 1'b0;
      sigmoid_table_488_0_sva <= 1'b0;
      sigmoid_table_488_5_sva <= 1'b0;
      sigmoid_table_487_0_sva <= 1'b0;
      sigmoid_table_486_0_sva <= 1'b0;
      sigmoid_table_485_0_sva <= 1'b0;
      sigmoid_table_485_2_sva <= 1'b0;
      sigmoid_table_485_4_sva <= 1'b0;
      sigmoid_table_484_0_sva <= 1'b0;
      sigmoid_table_484_4_sva <= 1'b0;
      sigmoid_table_483_0_sva <= 1'b0;
      sigmoid_table_482_1_sva <= 1'b0;
      sigmoid_table_482_3_sva <= 1'b0;
      sigmoid_table_480_1_sva <= 1'b0;
      sigmoid_table_479_8_sva <= 1'b0;
      sigmoid_table_478_8_sva <= 1'b0;
      sigmoid_table_477_8_sva <= 1'b0;
      sigmoid_table_476_8_sva <= 1'b0;
      sigmoid_table_475_8_sva <= 1'b0;
      sigmoid_table_474_8_sva <= 1'b0;
      sigmoid_table_473_3_sva <= 1'b0;
      sigmoid_table_473_8_sva <= 1'b0;
      sigmoid_table_472_0_sva <= 1'b0;
      sigmoid_table_472_2_sva <= 1'b0;
      sigmoid_table_472_8_sva <= 1'b0;
      sigmoid_table_471_0_sva <= 1'b0;
      sigmoid_table_471_8_sva <= 1'b0;
      sigmoid_table_470_0_sva <= 1'b0;
      sigmoid_table_470_6_sva <= 1'b0;
      sigmoid_table_470_8_sva <= 1'b0;
      sigmoid_table_469_1_sva <= 1'b0;
      sigmoid_table_469_6_sva <= 1'b0;
      sigmoid_table_469_8_sva <= 1'b0;
      sigmoid_table_468_4_sva <= 1'b0;
      sigmoid_table_468_6_sva <= 1'b0;
      sigmoid_table_468_8_sva <= 1'b0;
      sigmoid_table_467_4_sva <= 1'b0;
      sigmoid_table_467_6_sva <= 1'b0;
      sigmoid_table_467_8_sva <= 1'b0;
      sigmoid_table_466_6_sva <= 1'b0;
      sigmoid_table_466_8_sva <= 1'b0;
      sigmoid_table_465_6_sva <= 1'b0;
      sigmoid_table_465_8_sva <= 1'b0;
      sigmoid_table_464_3_sva <= 1'b0;
      sigmoid_table_464_6_sva <= 1'b0;
      sigmoid_table_464_8_sva <= 1'b0;
      sigmoid_table_463_0_sva <= 1'b0;
      sigmoid_table_463_2_sva <= 1'b0;
      sigmoid_table_463_6_sva <= 1'b0;
      sigmoid_table_463_8_sva <= 1'b0;
      sigmoid_table_462_0_sva <= 1'b0;
      sigmoid_table_462_6_sva <= 1'b0;
      sigmoid_table_462_8_sva <= 1'b0;
      sigmoid_table_461_8_sva <= 1'b0;
      sigmoid_table_460_1_sva <= 1'b0;
      sigmoid_table_460_8_sva <= 1'b0;
      sigmoid_table_459_8_sva <= 1'b0;
      sigmoid_table_458_8_sva <= 1'b0;
      sigmoid_table_457_8_sva <= 1'b0;
      sigmoid_table_456_0_sva <= 1'b0;
      sigmoid_table_456_5_sva <= 1'b0;
      sigmoid_table_456_8_sva <= 1'b0;
      sigmoid_table_455_0_sva <= 1'b0;
      sigmoid_table_455_3_sva <= 1'b0;
      sigmoid_table_455_5_sva <= 1'b0;
      sigmoid_table_455_8_sva <= 1'b0;
      sigmoid_table_454_5_sva <= 1'b0;
      sigmoid_table_454_8_sva <= 1'b0;
      sigmoid_table_453_5_sva <= 1'b0;
      sigmoid_table_453_8_sva <= 1'b0;
      sigmoid_table_452_5_sva <= 1'b0;
      sigmoid_table_452_8_sva <= 1'b0;
      sigmoid_table_451_8_sva <= 1'b0;
      sigmoid_table_450_0_sva <= 1'b0;
      sigmoid_table_450_8_sva <= 1'b0;
      sigmoid_table_449_4_sva <= 1'b0;
      sigmoid_table_449_8_sva <= 1'b0;
      sigmoid_table_448_4_sva <= 1'b0;
      sigmoid_table_448_8_sva <= 1'b0;
      sigmoid_table_447_4_sva <= 1'b0;
      sigmoid_table_447_8_sva <= 1'b0;
      sigmoid_table_446_0_sva <= 1'b0;
      sigmoid_table_446_8_sva <= 1'b0;
      sigmoid_table_445_1_sva <= 1'b0;
      sigmoid_table_445_3_sva <= 1'b0;
      sigmoid_table_445_8_sva <= 1'b0;
      sigmoid_table_444_8_sva <= 1'b0;
      sigmoid_table_443_8_sva <= 1'b0;
      sigmoid_table_442_8_sva <= 1'b0;
      sigmoid_table_441_0_sva <= 1'b0;
      sigmoid_table_440_1_sva <= 1'b0;
      sigmoid_table_438_0_sva <= 1'b0;
      sigmoid_table_438_2_sva <= 1'b0;
      sigmoid_table_437_1_sva <= 1'b0;
      sigmoid_table_434_0_sva <= 1'b0;
      sigmoid_table_434_3_sva <= 1'b0;
      sigmoid_table_432_2_sva <= 1'b0;
      sigmoid_table_431_0_sva <= 1'b0;
      sigmoid_table_428_0_sva <= 1'b0;
      sigmoid_table_427_4_sva <= 1'b0;
      sigmoid_table_426_4_sva <= 1'b0;
      sigmoid_table_425_0_sva <= 1'b0;
      sigmoid_table_425_4_sva <= 1'b0;
      sigmoid_table_422_0_sva <= 1'b0;
      sigmoid_table_422_3_sva <= 1'b0;
      sigmoid_table_420_2_sva <= 1'b0;
      sigmoid_table_419_1_sva <= 1'b0;
      sigmoid_table_418_7_sva <= 1'b0;
      sigmoid_table_417_0_sva <= 1'b0;
      sigmoid_table_417_7_sva <= 1'b0;
      sigmoid_table_416_1_sva <= 1'b0;
      sigmoid_table_416_7_sva <= 1'b0;
      sigmoid_table_415_7_sva <= 1'b0;
      sigmoid_table_414_7_sva <= 1'b0;
      sigmoid_table_413_7_sva <= 1'b0;
      sigmoid_table_412_0_sva <= 1'b0;
      sigmoid_table_412_7_sva <= 1'b0;
      sigmoid_table_411_5_sva <= 1'b0;
      sigmoid_table_411_7_sva <= 1'b0;
      sigmoid_table_410_5_sva <= 1'b0;
      sigmoid_table_410_7_sva <= 1'b0;
      sigmoid_table_409_1_sva <= 1'b0;
      sigmoid_table_409_3_sva <= 1'b0;
      sigmoid_table_409_5_sva <= 1'b0;
      sigmoid_table_409_7_sva <= 1'b0;
      sigmoid_table_408_3_sva <= 1'b0;
      sigmoid_table_408_5_sva <= 1'b0;
      sigmoid_table_408_7_sva <= 1'b0;
      sigmoid_table_407_5_sva <= 1'b0;
      sigmoid_table_407_7_sva <= 1'b0;
      sigmoid_table_406_2_sva <= 1'b0;
      sigmoid_table_406_5_sva <= 1'b0;
      sigmoid_table_406_7_sva <= 1'b0;
      sigmoid_table_405_0_sva <= 1'b0;
      sigmoid_table_405_5_sva <= 1'b0;
      sigmoid_table_405_7_sva <= 1'b0;
      sigmoid_table_404_7_sva <= 1'b0;
      sigmoid_table_403_0_sva <= 1'b0;
      sigmoid_table_403_7_sva <= 1'b0;
      sigmoid_table_402_7_sva <= 1'b0;
      sigmoid_table_401_0_sva <= 1'b0;
      sigmoid_table_401_7_sva <= 1'b0;
      sigmoid_table_400_4_sva <= 1'b0;
      sigmoid_table_400_7_sva <= 1'b0;
      sigmoid_table_399_0_sva <= 1'b0;
      sigmoid_table_399_2_sva <= 1'b0;
      sigmoid_table_399_4_sva <= 1'b0;
      sigmoid_table_399_7_sva <= 1'b0;
      sigmoid_table_398_4_sva <= 1'b0;
      sigmoid_table_398_7_sva <= 1'b0;
      sigmoid_table_397_0_sva <= 1'b0;
      sigmoid_table_397_4_sva <= 1'b0;
      sigmoid_table_397_7_sva <= 1'b0;
      sigmoid_table_396_7_sva <= 1'b0;
      sigmoid_table_395_0_sva <= 1'b0;
      sigmoid_table_395_7_sva <= 1'b0;
      sigmoid_table_394_3_sva <= 1'b0;
      sigmoid_table_394_7_sva <= 1'b0;
      sigmoid_table_393_1_sva <= 1'b0;
      sigmoid_table_393_3_sva <= 1'b0;
      sigmoid_table_393_7_sva <= 1'b0;
      sigmoid_table_392_3_sva <= 1'b0;
      sigmoid_table_392_7_sva <= 1'b0;
      sigmoid_table_391_7_sva <= 1'b0;
      sigmoid_table_390_2_sva <= 1'b0;
      sigmoid_table_390_7_sva <= 1'b0;
      sigmoid_table_389_1_sva <= 1'b0;
      sigmoid_table_389_7_sva <= 1'b0;
      sigmoid_table_388_7_sva <= 1'b0;
      sigmoid_table_386_0_sva <= 1'b0;
      sigmoid_table_384_1_sva <= 1'b0;
      sigmoid_table_381_0_sva <= 1'b0;
      sigmoid_table_381_2_sva <= 1'b0;
      sigmoid_table_379_0_sva <= 1'b0;
      sigmoid_table_376_0_sva <= 1'b0;
      sigmoid_table_375_3_sva <= 1'b0;
      sigmoid_table_374_1_sva <= 1'b0;
      sigmoid_table_374_3_sva <= 1'b0;
      sigmoid_table_373_3_sva <= 1'b0;
      sigmoid_table_371_0_sva <= 1'b0;
      sigmoid_table_371_2_sva <= 1'b0;
      sigmoid_table_370_2_sva <= 1'b0;
      sigmoid_table_368_0_sva <= 1'b0;
      sigmoid_table_366_6_sva <= 1'b0;
      sigmoid_table_365_0_sva <= 1'b0;
      sigmoid_table_365_6_sva <= 1'b0;
      sigmoid_table_364_6_sva <= 1'b0;
      sigmoid_table_363_1_sva <= 1'b0;
      sigmoid_table_363_6_sva <= 1'b0;
      sigmoid_table_362_0_sva <= 1'b0;
      sigmoid_table_362_6_sva <= 1'b0;
      sigmoid_table_361_6_sva <= 1'b0;
      sigmoid_table_360_4_sva <= 1'b0;
      sigmoid_table_360_6_sva <= 1'b0;
      sigmoid_table_359_0_sva <= 1'b0;
      sigmoid_table_359_2_sva <= 1'b0;
      sigmoid_table_359_4_sva <= 1'b0;
      sigmoid_table_359_6_sva <= 1'b0;
      sigmoid_table_358_2_sva <= 1'b0;
      sigmoid_table_358_4_sva <= 1'b0;
      sigmoid_table_358_6_sva <= 1'b0;
      sigmoid_table_357_4_sva <= 1'b0;
      sigmoid_table_357_6_sva <= 1'b0;
      sigmoid_table_356_1_sva <= 1'b0;
      sigmoid_table_356_4_sva <= 1'b0;
      sigmoid_table_356_6_sva <= 1'b0;
      sigmoid_table_355_0_sva <= 1'b0;
      sigmoid_table_355_4_sva <= 1'b0;
      sigmoid_table_355_6_sva <= 1'b0;
      sigmoid_table_354_6_sva <= 1'b0;
      sigmoid_table_353_6_sva <= 1'b0;
      sigmoid_table_352_0_sva <= 1'b0;
      sigmoid_table_352_6_sva <= 1'b0;
      sigmoid_table_351_6_sva <= 1'b0;
      sigmoid_table_350_3_sva <= 1'b0;
      sigmoid_table_350_6_sva <= 1'b0;
      sigmoid_table_349_1_sva <= 1'b0;
      sigmoid_table_349_3_sva <= 1'b0;
      sigmoid_table_349_6_sva <= 1'b0;
      sigmoid_table_348_0_sva <= 1'b0;
      sigmoid_table_348_3_sva <= 1'b0;
      sigmoid_table_348_6_sva <= 1'b0;
      sigmoid_table_347_3_sva <= 1'b0;
      sigmoid_table_347_6_sva <= 1'b0;
      sigmoid_table_346_6_sva <= 1'b0;
      sigmoid_table_345_6_sva <= 1'b0;
      sigmoid_table_344_0_sva <= 1'b0;
      sigmoid_table_344_2_sva <= 1'b0;
      sigmoid_table_344_6_sva <= 1'b0;
      sigmoid_table_343_2_sva <= 1'b0;
      sigmoid_table_343_6_sva <= 1'b0;
      sigmoid_table_342_6_sva <= 1'b0;
      sigmoid_table_341_1_sva <= 1'b0;
      sigmoid_table_341_6_sva <= 1'b0;
      sigmoid_table_340_0_sva <= 1'b0;
      sigmoid_table_340_6_sva <= 1'b0;
      sigmoid_table_339_6_sva <= 1'b0;
      sigmoid_table_336_0_sva <= 1'b0;
      sigmoid_table_333_1_sva <= 1'b0;
      sigmoid_table_332_1_sva <= 1'b0;
      sigmoid_table_331_0_sva <= 1'b0;
      sigmoid_table_327_0_sva <= 1'b0;
      sigmoid_table_327_2_sva <= 1'b0;
      sigmoid_table_326_0_sva <= 1'b0;
      sigmoid_table_326_2_sva <= 1'b0;
      sigmoid_table_325_2_sva <= 1'b0;
      sigmoid_table_323_1_sva <= 1'b0;
      sigmoid_table_322_1_sva <= 1'b0;
      sigmoid_table_321_0_sva <= 1'b0;
      sigmoid_table_319_5_sva <= 1'b0;
      sigmoid_table_318_5_sva <= 1'b0;
      sigmoid_table_317_5_sva <= 1'b0;
      sigmoid_table_316_0_sva <= 1'b0;
      sigmoid_table_316_5_sva <= 1'b0;
      sigmoid_table_315_0_sva <= 1'b0;
      sigmoid_table_315_5_sva <= 1'b0;
      sigmoid_table_314_5_sva <= 1'b0;
      sigmoid_table_313_3_sva <= 1'b0;
      sigmoid_table_313_5_sva <= 1'b0;
      sigmoid_table_312_3_sva <= 1'b0;
      sigmoid_table_312_5_sva <= 1'b0;
      sigmoid_table_311_1_sva <= 1'b0;
      sigmoid_table_311_3_sva <= 1'b0;
      sigmoid_table_311_5_sva <= 1'b0;
      sigmoid_table_310_0_sva <= 1'b0;
      sigmoid_table_310_3_sva <= 1'b0;
      sigmoid_table_310_5_sva <= 1'b0;
      sigmoid_table_309_0_sva <= 1'b0;
      sigmoid_table_309_3_sva <= 1'b0;
      sigmoid_table_309_5_sva <= 1'b0;
      sigmoid_table_308_3_sva <= 1'b0;
      sigmoid_table_308_5_sva <= 1'b0;
      sigmoid_table_307_5_sva <= 1'b0;
      sigmoid_table_306_5_sva <= 1'b0;
      sigmoid_table_305_5_sva <= 1'b0;
      sigmoid_table_304_5_sva <= 1'b0;
      sigmoid_table_303_0_sva <= 1'b0;
      sigmoid_table_303_2_sva <= 1'b0;
      sigmoid_table_303_5_sva <= 1'b0;
      sigmoid_table_302_0_sva <= 1'b0;
      sigmoid_table_302_2_sva <= 1'b0;
      sigmoid_table_302_5_sva <= 1'b0;
      sigmoid_table_301_2_sva <= 1'b0;
      sigmoid_table_301_5_sva <= 1'b0;
      sigmoid_table_300_5_sva <= 1'b0;
      sigmoid_table_299_5_sva <= 1'b0;
      sigmoid_table_298_1_sva <= 1'b0;
      sigmoid_table_298_5_sva <= 1'b0;
      sigmoid_table_297_1_sva <= 1'b0;
      sigmoid_table_297_5_sva <= 1'b0;
      sigmoid_table_296_0_sva <= 1'b0;
      sigmoid_table_296_5_sva <= 1'b0;
      sigmoid_table_295_0_sva <= 1'b0;
      sigmoid_table_295_5_sva <= 1'b0;
      sigmoid_table_294_5_sva <= 1'b0;
      sigmoid_table_293_5_sva <= 1'b0;
      sigmoid_table_287_0_sva <= 1'b0;
      sigmoid_table_286_0_sva <= 1'b0;
      sigmoid_table_281_1_sva <= 1'b0;
      sigmoid_table_280_1_sva <= 1'b0;
      sigmoid_table_279_1_sva <= 1'b0;
      sigmoid_table_278_0_sva <= 1'b0;
      sigmoid_table_277_0_sva <= 1'b0;
      sigmoid_table_276_0_sva <= 1'b0;
      sigmoid_table_273_4_sva <= 1'b0;
      sigmoid_table_272_4_sva <= 1'b0;
      sigmoid_table_271_4_sva <= 1'b0;
      sigmoid_table_270_4_sva <= 1'b0;
      sigmoid_table_269_4_sva <= 1'b0;
      sigmoid_table_268_4_sva <= 1'b0;
      sigmoid_table_267_0_sva <= 1'b0;
      sigmoid_table_267_2_sva <= 1'b0;
      sigmoid_table_267_4_sva <= 1'b0;
      sigmoid_table_266_0_sva <= 1'b0;
      sigmoid_table_266_2_sva <= 1'b0;
      sigmoid_table_266_4_sva <= 1'b0;
      sigmoid_table_265_0_sva <= 1'b0;
      sigmoid_table_265_2_sva <= 1'b0;
      sigmoid_table_265_4_sva <= 1'b0;
      sigmoid_table_264_2_sva <= 1'b0;
      sigmoid_table_264_4_sva <= 1'b0;
      sigmoid_table_263_2_sva <= 1'b0;
      sigmoid_table_263_4_sva <= 1'b0;
      sigmoid_table_262_2_sva <= 1'b0;
      sigmoid_table_262_4_sva <= 1'b0;
      sigmoid_table_261_4_sva <= 1'b0;
      sigmoid_table_260_4_sva <= 1'b0;
      sigmoid_table_259_4_sva <= 1'b0;
      sigmoid_table_258_1_sva <= 1'b0;
      sigmoid_table_258_4_sva <= 1'b0;
      sigmoid_table_257_1_sva <= 1'b0;
      sigmoid_table_257_4_sva <= 1'b0;
      sigmoid_table_256_1_sva <= 1'b0;
      sigmoid_table_256_4_sva <= 1'b0;
      sigmoid_table_255_1_sva <= 1'b0;
      sigmoid_table_255_4_sva <= 1'b0;
      sigmoid_table_254_0_sva <= 1'b0;
      sigmoid_table_254_4_sva <= 1'b0;
      sigmoid_table_253_0_sva <= 1'b0;
      sigmoid_table_253_4_sva <= 1'b0;
      sigmoid_table_252_0_sva <= 1'b0;
      sigmoid_table_252_4_sva <= 1'b0;
      sigmoid_table_251_0_sva <= 1'b0;
      sigmoid_table_251_4_sva <= 1'b0;
      sigmoid_table_250_4_sva <= 1'b0;
      sigmoid_table_249_4_sva <= 1'b0;
      sigmoid_table_248_4_sva <= 1'b0;
      sigmoid_table_247_4_sva <= 1'b0;
      sigmoid_table_238_0_sva <= 1'b0;
      sigmoid_table_237_0_sva <= 1'b0;
      sigmoid_table_236_0_sva <= 1'b0;
      sigmoid_table_235_0_sva <= 1'b0;
      sigmoid_table_234_0_sva <= 1'b0;
      sigmoid_table_228_3_sva <= 1'b0;
      sigmoid_table_227_3_sva <= 1'b0;
      sigmoid_table_226_3_sva <= 1'b0;
      sigmoid_table_225_3_sva <= 1'b0;
      sigmoid_table_224_3_sva <= 1'b0;
      sigmoid_table_223_3_sva <= 1'b0;
      sigmoid_table_222_1_sva <= 1'b0;
      sigmoid_table_222_3_sva <= 1'b0;
      sigmoid_table_221_1_sva <= 1'b0;
      sigmoid_table_221_3_sva <= 1'b0;
      sigmoid_table_220_1_sva <= 1'b0;
      sigmoid_table_220_3_sva <= 1'b0;
      sigmoid_table_219_1_sva <= 1'b0;
      sigmoid_table_219_3_sva <= 1'b0;
      sigmoid_table_218_1_sva <= 1'b0;
      sigmoid_table_218_3_sva <= 1'b0;
      sigmoid_table_217_1_sva <= 1'b0;
      sigmoid_table_217_3_sva <= 1'b0;
      sigmoid_table_216_0_sva <= 1'b0;
      sigmoid_table_216_3_sva <= 1'b0;
      sigmoid_table_215_0_sva <= 1'b0;
      sigmoid_table_215_3_sva <= 1'b0;
      sigmoid_table_214_0_sva <= 1'b0;
      sigmoid_table_214_3_sva <= 1'b0;
      sigmoid_table_213_0_sva <= 1'b0;
      sigmoid_table_213_3_sva <= 1'b0;
      sigmoid_table_212_0_sva <= 1'b0;
      sigmoid_table_212_3_sva <= 1'b0;
      sigmoid_table_211_0_sva <= 1'b0;
      sigmoid_table_211_3_sva <= 1'b0;
      sigmoid_table_210_0_sva <= 1'b0;
      sigmoid_table_210_3_sva <= 1'b0;
      sigmoid_table_209_3_sva <= 1'b0;
      sigmoid_table_208_3_sva <= 1'b0;
      sigmoid_table_207_3_sva <= 1'b0;
      sigmoid_table_206_3_sva <= 1'b0;
      sigmoid_table_205_3_sva <= 1'b0;
      sigmoid_table_204_3_sva <= 1'b0;
      sigmoid_table_203_3_sva <= 1'b0;
      sigmoid_table_202_3_sva <= 1'b0;
      sigmoid_table_183_0_sva <= 1'b0;
      sigmoid_table_183_2_sva <= 1'b0;
      sigmoid_table_182_0_sva <= 1'b0;
      sigmoid_table_182_2_sva <= 1'b0;
      sigmoid_table_181_0_sva <= 1'b0;
      sigmoid_table_181_2_sva <= 1'b0;
      sigmoid_table_180_0_sva <= 1'b0;
      sigmoid_table_180_2_sva <= 1'b0;
      sigmoid_table_179_0_sva <= 1'b0;
      sigmoid_table_179_2_sva <= 1'b0;
      sigmoid_table_178_0_sva <= 1'b0;
      sigmoid_table_178_2_sva <= 1'b0;
      sigmoid_table_177_0_sva <= 1'b0;
      sigmoid_table_177_2_sva <= 1'b0;
      sigmoid_table_176_0_sva <= 1'b0;
      sigmoid_table_176_2_sva <= 1'b0;
      sigmoid_table_175_0_sva <= 1'b0;
      sigmoid_table_175_2_sva <= 1'b0;
      sigmoid_table_174_0_sva <= 1'b0;
      sigmoid_table_174_2_sva <= 1'b0;
      sigmoid_table_173_0_sva <= 1'b0;
      sigmoid_table_173_2_sva <= 1'b0;
      sigmoid_table_172_0_sva <= 1'b0;
      sigmoid_table_172_2_sva <= 1'b0;
      sigmoid_table_171_2_sva <= 1'b0;
      sigmoid_table_170_2_sva <= 1'b0;
      sigmoid_table_169_2_sva <= 1'b0;
      sigmoid_table_168_2_sva <= 1'b0;
      sigmoid_table_167_2_sva <= 1'b0;
      sigmoid_table_166_2_sva <= 1'b0;
      sigmoid_table_165_2_sva <= 1'b0;
      sigmoid_table_164_2_sva <= 1'b0;
      sigmoid_table_163_2_sva <= 1'b0;
      sigmoid_table_162_2_sva <= 1'b0;
      sigmoid_table_161_2_sva <= 1'b0;
      sigmoid_table_160_2_sva <= 1'b0;
      sigmoid_table_159_2_sva <= 1'b0;
      sigmoid_table_158_2_sva <= 1'b0;
      sigmoid_table_138_1_sva <= 1'b0;
      sigmoid_table_137_1_sva <= 1'b0;
      sigmoid_table_136_1_sva <= 1'b0;
      sigmoid_table_135_1_sva <= 1'b0;
      sigmoid_table_134_1_sva <= 1'b0;
      sigmoid_table_133_1_sva <= 1'b0;
      sigmoid_table_132_1_sva <= 1'b0;
      sigmoid_table_131_1_sva <= 1'b0;
      sigmoid_table_130_1_sva <= 1'b0;
      sigmoid_table_129_1_sva <= 1'b0;
      sigmoid_table_128_1_sva <= 1'b0;
      sigmoid_table_127_1_sva <= 1'b0;
      sigmoid_table_126_1_sva <= 1'b0;
      sigmoid_table_125_1_sva <= 1'b0;
      sigmoid_table_124_1_sva <= 1'b0;
      sigmoid_table_123_1_sva <= 1'b0;
      sigmoid_table_122_1_sva <= 1'b0;
      sigmoid_table_121_1_sva <= 1'b0;
      sigmoid_table_120_1_sva <= 1'b0;
      sigmoid_table_119_1_sva <= 1'b0;
      sigmoid_table_118_1_sva <= 1'b0;
      sigmoid_table_117_1_sva <= 1'b0;
      sigmoid_table_116_1_sva <= 1'b0;
      sigmoid_table_115_1_sva <= 1'b0;
      sigmoid_table_114_1_sva <= 1'b0;
      sigmoid_table_113_1_sva <= 1'b0;
      sigmoid_table_112_0_sva <= 1'b0;
      sigmoid_table_111_0_sva <= 1'b0;
      sigmoid_table_110_0_sva <= 1'b0;
      sigmoid_table_109_0_sva <= 1'b0;
      sigmoid_table_108_0_sva <= 1'b0;
      sigmoid_table_107_0_sva <= 1'b0;
      sigmoid_table_106_0_sva <= 1'b0;
      sigmoid_table_105_0_sva <= 1'b0;
      sigmoid_table_104_0_sva <= 1'b0;
      sigmoid_table_103_0_sva <= 1'b0;
      sigmoid_table_102_0_sva <= 1'b0;
      sigmoid_table_101_0_sva <= 1'b0;
      sigmoid_table_100_0_sva <= 1'b0;
      sigmoid_table_99_0_sva <= 1'b0;
      sigmoid_table_98_0_sva <= 1'b0;
      sigmoid_table_97_0_sva <= 1'b0;
      sigmoid_table_96_0_sva <= 1'b0;
      sigmoid_table_95_0_sva <= 1'b0;
      sigmoid_table_94_0_sva <= 1'b0;
      sigmoid_table_93_0_sva <= 1'b0;
      sigmoid_table_92_0_sva <= 1'b0;
      sigmoid_table_91_0_sva <= 1'b0;
      sigmoid_table_90_0_sva <= 1'b0;
      sigmoid_table_89_0_sva <= 1'b0;
      sigmoid_table_88_0_sva <= 1'b0;
      sigmoid_table_87_0_sva <= 1'b0;
      sigmoid_table_86_0_sva <= 1'b0;
      sigmoid_table_85_0_sva <= 1'b0;
      sigmoid_table_84_0_sva <= 1'b0;
      sigmoid_table_83_0_sva <= 1'b0;
      sigmoid_table_82_0_sva <= 1'b0;
      sigmoid_table_81_0_sva <= 1'b0;
      sigmoid_table_80_0_sva <= 1'b0;
      sigmoid_table_79_0_sva <= 1'b0;
      sigmoid_table_78_0_sva <= 1'b0;
      sigmoid_table_77_0_sva <= 1'b0;
      sigmoid_table_76_0_sva <= 1'b0;
      sigmoid_table_75_0_sva <= 1'b0;
      sigmoid_table_74_0_sva <= 1'b0;
      sigmoid_table_73_0_sva <= 1'b0;
      sigmoid_table_72_0_sva <= 1'b0;
      sigmoid_table_71_0_sva <= 1'b0;
      sigmoid_table_70_0_sva <= 1'b0;
      sigmoid_table_69_0_sva <= 1'b0;
    end
    else if ( sigmoid_table_and_cse ) begin
      sigmoid_table_1023_0_sva <= sigmoid_table_1023_0_sva_dfm_1;
      sigmoid_table_1022_0_sva <= sigmoid_table_1022_0_sva_dfm_1;
      sigmoid_table_1021_0_sva <= sigmoid_table_1021_0_sva_dfm_1;
      sigmoid_table_1020_0_sva <= sigmoid_table_1020_0_sva_dfm_1;
      sigmoid_table_1019_0_sva <= sigmoid_table_1019_0_sva_dfm_1;
      sigmoid_table_1018_0_sva <= sigmoid_table_1018_0_sva_dfm_1;
      sigmoid_table_1017_0_sva <= sigmoid_table_1017_0_sva_dfm_1;
      sigmoid_table_1016_0_sva <= sigmoid_table_1016_0_sva_dfm_1;
      sigmoid_table_1015_0_sva <= sigmoid_table_1015_0_sva_dfm_1;
      sigmoid_table_1014_0_sva <= sigmoid_table_1014_0_sva_dfm_1;
      sigmoid_table_1013_0_sva <= sigmoid_table_1013_0_sva_dfm_1;
      sigmoid_table_1012_0_sva <= sigmoid_table_1012_0_sva_dfm_1;
      sigmoid_table_1011_0_sva <= sigmoid_table_1011_0_sva_dfm_1;
      sigmoid_table_1010_0_sva <= sigmoid_table_1010_0_sva_dfm_1;
      sigmoid_table_1009_0_sva <= sigmoid_table_1009_0_sva_dfm_1;
      sigmoid_table_1008_0_sva <= sigmoid_table_1008_0_sva_dfm_1;
      sigmoid_table_1007_0_sva <= sigmoid_table_1007_0_sva_dfm_1;
      sigmoid_table_1006_0_sva <= sigmoid_table_1006_0_sva_dfm_1;
      sigmoid_table_1005_0_sva <= sigmoid_table_1005_0_sva_dfm_1;
      sigmoid_table_1004_0_sva <= sigmoid_table_1004_0_sva_dfm_1;
      sigmoid_table_1003_0_sva <= sigmoid_table_1003_0_sva_dfm_1;
      sigmoid_table_1002_0_sva <= sigmoid_table_1002_0_sva_dfm_1;
      sigmoid_table_1001_0_sva <= sigmoid_table_1001_0_sva_dfm_1;
      sigmoid_table_1000_0_sva <= sigmoid_table_1000_0_sva_dfm_1;
      sigmoid_table_999_0_sva <= sigmoid_table_999_0_sva_dfm_1;
      sigmoid_table_998_0_sva <= sigmoid_table_998_0_sva_dfm_1;
      sigmoid_table_997_0_sva <= sigmoid_table_997_0_sva_dfm_1;
      sigmoid_table_996_0_sva <= sigmoid_table_996_0_sva_dfm_1;
      sigmoid_table_995_0_sva <= sigmoid_table_995_0_sva_dfm_1;
      sigmoid_table_994_0_sva <= sigmoid_table_994_0_sva_dfm_1;
      sigmoid_table_993_0_sva <= sigmoid_table_993_0_sva_dfm_1;
      sigmoid_table_992_0_sva <= sigmoid_table_992_0_sva_dfm_1;
      sigmoid_table_991_0_sva <= sigmoid_table_991_0_sva_dfm_1;
      sigmoid_table_990_0_sva <= sigmoid_table_990_0_sva_dfm_1;
      sigmoid_table_989_0_sva <= sigmoid_table_989_0_sva_dfm_1;
      sigmoid_table_988_0_sva <= sigmoid_table_988_0_sva_dfm_1;
      sigmoid_table_987_0_sva <= sigmoid_table_987_0_sva_dfm_1;
      sigmoid_table_986_0_sva <= sigmoid_table_986_0_sva_dfm_1;
      sigmoid_table_985_0_sva <= sigmoid_table_985_0_sva_dfm_1;
      sigmoid_table_984_0_sva <= sigmoid_table_984_0_sva_dfm_1;
      sigmoid_table_983_0_sva <= sigmoid_table_983_0_sva_dfm_1;
      sigmoid_table_982_0_sva <= sigmoid_table_982_0_sva_dfm_1;
      sigmoid_table_981_0_sva <= sigmoid_table_981_0_sva_dfm_1;
      sigmoid_table_980_0_sva <= sigmoid_table_980_0_sva_dfm_1;
      sigmoid_table_979_0_sva <= sigmoid_table_979_0_sva_dfm_1;
      sigmoid_table_978_0_sva <= sigmoid_table_978_0_sva_dfm_1;
      sigmoid_table_977_0_sva <= sigmoid_table_977_0_sva_dfm_1;
      sigmoid_table_976_0_sva <= sigmoid_table_976_0_sva_dfm_1;
      sigmoid_table_975_0_sva <= sigmoid_table_975_0_sva_dfm_1;
      sigmoid_table_974_0_sva <= sigmoid_table_974_0_sva_dfm_1;
      sigmoid_table_973_0_sva <= sigmoid_table_973_0_sva_dfm_1;
      sigmoid_table_972_0_sva <= sigmoid_table_972_0_sva_dfm_1;
      sigmoid_table_971_0_sva <= sigmoid_table_971_0_sva_dfm_1;
      sigmoid_table_970_0_sva <= sigmoid_table_970_0_sva_dfm_1;
      sigmoid_table_969_0_sva <= sigmoid_table_969_0_sva_dfm_1;
      sigmoid_table_968_0_sva <= sigmoid_table_968_0_sva_dfm_1;
      sigmoid_table_967_0_sva <= sigmoid_table_967_0_sva_dfm_1;
      sigmoid_table_966_0_sva <= sigmoid_table_966_0_sva_dfm_1;
      sigmoid_table_965_0_sva <= sigmoid_table_965_0_sva_dfm_1;
      sigmoid_table_964_0_sva <= sigmoid_table_964_0_sva_dfm_1;
      sigmoid_table_963_0_sva <= sigmoid_table_963_0_sva_dfm_1;
      sigmoid_table_962_0_sva <= sigmoid_table_962_0_sva_dfm_1;
      sigmoid_table_961_0_sva <= sigmoid_table_961_0_sva_dfm_1;
      sigmoid_table_960_0_sva <= sigmoid_table_960_0_sva_dfm_1;
      sigmoid_table_959_0_sva <= sigmoid_table_959_0_sva_dfm_1;
      sigmoid_table_958_0_sva <= sigmoid_table_958_0_sva_dfm_1;
      sigmoid_table_957_0_sva <= sigmoid_table_957_0_sva_dfm_1;
      sigmoid_table_956_0_sva <= sigmoid_table_956_0_sva_dfm_1;
      sigmoid_table_955_0_sva <= sigmoid_table_955_0_sva_dfm_1;
      sigmoid_table_954_1_sva <= sigmoid_table_954_1_sva_dfm_1;
      sigmoid_table_953_1_sva <= sigmoid_table_953_1_sva_dfm_1;
      sigmoid_table_952_1_sva <= sigmoid_table_952_1_sva_dfm_1;
      sigmoid_table_951_1_sva <= sigmoid_table_951_1_sva_dfm_1;
      sigmoid_table_950_1_sva <= sigmoid_table_950_1_sva_dfm_1;
      sigmoid_table_949_1_sva <= sigmoid_table_949_1_sva_dfm_1;
      sigmoid_table_948_1_sva <= sigmoid_table_948_1_sva_dfm_1;
      sigmoid_table_947_1_sva <= sigmoid_table_947_1_sva_dfm_1;
      sigmoid_table_946_1_sva <= sigmoid_table_946_1_sva_dfm_1;
      sigmoid_table_945_1_sva <= sigmoid_table_945_1_sva_dfm_1;
      sigmoid_table_944_1_sva <= sigmoid_table_944_1_sva_dfm_1;
      sigmoid_table_943_1_sva <= sigmoid_table_943_1_sva_dfm_1;
      sigmoid_table_942_1_sva <= sigmoid_table_942_1_sva_dfm_1;
      sigmoid_table_941_1_sva <= sigmoid_table_941_1_sva_dfm_1;
      sigmoid_table_940_1_sva <= sigmoid_table_940_1_sva_dfm_1;
      sigmoid_table_939_1_sva <= sigmoid_table_939_1_sva_dfm_1;
      sigmoid_table_938_1_sva <= sigmoid_table_938_1_sva_dfm_1;
      sigmoid_table_937_1_sva <= sigmoid_table_937_1_sva_dfm_1;
      sigmoid_table_936_1_sva <= sigmoid_table_936_1_sva_dfm_1;
      sigmoid_table_935_1_sva <= sigmoid_table_935_1_sva_dfm_1;
      sigmoid_table_934_1_sva <= sigmoid_table_934_1_sva_dfm_1;
      sigmoid_table_933_1_sva <= sigmoid_table_933_1_sva_dfm_1;
      sigmoid_table_932_1_sva <= sigmoid_table_932_1_sva_dfm_1;
      sigmoid_table_931_1_sva <= sigmoid_table_931_1_sva_dfm_1;
      sigmoid_table_930_1_sva <= sigmoid_table_930_1_sva_dfm_1;
      sigmoid_table_929_1_sva <= sigmoid_table_929_1_sva_dfm_1;
      sigmoid_table_928_1_sva <= sigmoid_table_928_1_sva_dfm_1;
      sigmoid_table_927_1_sva <= sigmoid_table_927_1_sva_dfm_1;
      sigmoid_table_926_1_sva <= sigmoid_table_926_1_sva_dfm_1;
      sigmoid_table_925_1_sva <= sigmoid_table_925_1_sva_dfm_1;
      sigmoid_table_924_1_sva <= sigmoid_table_924_1_sva_dfm_1;
      sigmoid_table_923_1_sva <= sigmoid_table_923_1_sva_dfm_1;
      sigmoid_table_922_1_sva <= sigmoid_table_922_1_sva_dfm_1;
      sigmoid_table_921_1_sva <= sigmoid_table_921_1_sva_dfm_1;
      sigmoid_table_920_1_sva <= sigmoid_table_920_1_sva_dfm_1;
      sigmoid_table_919_1_sva <= sigmoid_table_919_1_sva_dfm_1;
      sigmoid_table_918_1_sva <= sigmoid_table_918_1_sva_dfm_1;
      sigmoid_table_917_1_sva <= sigmoid_table_917_1_sva_dfm_1;
      sigmoid_table_916_1_sva <= sigmoid_table_916_1_sva_dfm_1;
      sigmoid_table_915_1_sva <= sigmoid_table_915_1_sva_dfm_1;
      sigmoid_table_914_1_sva <= sigmoid_table_914_1_sva_dfm_1;
      sigmoid_table_913_1_sva <= sigmoid_table_913_1_sva_dfm_1;
      sigmoid_table_912_1_sva <= sigmoid_table_912_1_sva_dfm_1;
      sigmoid_table_911_1_sva <= sigmoid_table_911_1_sva_dfm_1;
      sigmoid_table_910_2_sva <= sigmoid_table_910_2_sva_dfm_1;
      sigmoid_table_909_2_sva <= sigmoid_table_909_2_sva_dfm_1;
      sigmoid_table_908_2_sva <= sigmoid_table_908_2_sva_dfm_1;
      sigmoid_table_907_2_sva <= sigmoid_table_907_2_sva_dfm_1;
      sigmoid_table_906_2_sva <= sigmoid_table_906_2_sva_dfm_1;
      sigmoid_table_905_2_sva <= sigmoid_table_905_2_sva_dfm_1;
      sigmoid_table_904_2_sva <= sigmoid_table_904_2_sva_dfm_1;
      sigmoid_table_903_2_sva <= sigmoid_table_903_2_sva_dfm_1;
      sigmoid_table_902_2_sva <= sigmoid_table_902_2_sva_dfm_1;
      sigmoid_table_901_2_sva <= sigmoid_table_901_2_sva_dfm_1;
      sigmoid_table_900_2_sva <= sigmoid_table_900_2_sva_dfm_1;
      sigmoid_table_899_2_sva <= sigmoid_table_899_2_sva_dfm_1;
      sigmoid_table_898_2_sva <= sigmoid_table_898_2_sva_dfm_1;
      sigmoid_table_897_2_sva <= sigmoid_table_897_2_sva_dfm_1;
      sigmoid_table_896_2_sva <= sigmoid_table_896_2_sva_dfm_1;
      sigmoid_table_895_2_sva <= sigmoid_table_895_2_sva_dfm_1;
      sigmoid_table_894_2_sva <= sigmoid_table_894_2_sva_dfm_1;
      sigmoid_table_893_2_sva <= sigmoid_table_893_2_sva_dfm_1;
      sigmoid_table_892_2_sva <= sigmoid_table_892_2_sva_dfm_1;
      sigmoid_table_891_2_sva <= sigmoid_table_891_2_sva_dfm_1;
      sigmoid_table_890_2_sva <= sigmoid_table_890_2_sva_dfm_1;
      sigmoid_table_889_2_sva <= sigmoid_table_889_2_sva_dfm_1;
      sigmoid_table_888_2_sva <= sigmoid_table_888_2_sva_dfm_1;
      sigmoid_table_887_2_sva <= sigmoid_table_887_2_sva_dfm_1;
      sigmoid_table_886_2_sva <= sigmoid_table_886_2_sva_dfm_1;
      sigmoid_table_885_2_sva <= sigmoid_table_885_2_sva_dfm_1;
      sigmoid_table_884_2_sva <= sigmoid_table_884_2_sva_dfm_1;
      sigmoid_table_883_2_sva <= sigmoid_table_883_2_sva_dfm_1;
      sigmoid_table_882_2_sva <= sigmoid_table_882_2_sva_dfm_1;
      sigmoid_table_881_2_sva <= sigmoid_table_881_2_sva_dfm_1;
      sigmoid_table_880_2_sva <= sigmoid_table_880_2_sva_dfm_1;
      sigmoid_table_879_2_sva <= sigmoid_table_879_2_sva_dfm_1;
      sigmoid_table_878_2_sva <= sigmoid_table_878_2_sva_dfm_1;
      sigmoid_table_877_2_sva <= sigmoid_table_877_2_sva_dfm_1;
      sigmoid_table_876_2_sva <= sigmoid_table_876_2_sva_dfm_1;
      sigmoid_table_875_2_sva <= sigmoid_table_875_2_sva_dfm_1;
      sigmoid_table_874_2_sva <= sigmoid_table_874_2_sva_dfm_1;
      sigmoid_table_873_2_sva <= sigmoid_table_873_2_sva_dfm_1;
      sigmoid_table_872_2_sva <= sigmoid_table_872_2_sva_dfm_1;
      sigmoid_table_871_2_sva <= sigmoid_table_871_2_sva_dfm_1;
      sigmoid_table_870_2_sva <= sigmoid_table_870_2_sva_dfm_1;
      sigmoid_table_869_2_sva <= sigmoid_table_869_2_sva_dfm_1;
      sigmoid_table_868_2_sva <= sigmoid_table_868_2_sva_dfm_1;
      sigmoid_table_867_2_sva <= sigmoid_table_867_2_sva_dfm_1;
      sigmoid_table_866_0_sva <= sigmoid_table_866_0_sva_dfm_1;
      sigmoid_table_866_3_sva <= sigmoid_table_866_3_sva_dfm_1;
      sigmoid_table_865_0_sva <= sigmoid_table_865_0_sva_dfm_1;
      sigmoid_table_865_3_sva <= sigmoid_table_865_3_sva_dfm_1;
      sigmoid_table_864_0_sva <= sigmoid_table_864_0_sva_dfm_1;
      sigmoid_table_864_3_sva <= sigmoid_table_864_3_sva_dfm_1;
      sigmoid_table_863_0_sva <= sigmoid_table_863_0_sva_dfm_1;
      sigmoid_table_863_3_sva <= sigmoid_table_863_3_sva_dfm_1;
      sigmoid_table_862_0_sva <= sigmoid_table_862_0_sva_dfm_1;
      sigmoid_table_862_3_sva <= sigmoid_table_862_3_sva_dfm_1;
      sigmoid_table_861_0_sva <= sigmoid_table_861_0_sva_dfm_1;
      sigmoid_table_861_3_sva <= sigmoid_table_861_3_sva_dfm_1;
      sigmoid_table_860_0_sva <= sigmoid_table_860_0_sva_dfm_1;
      sigmoid_table_860_3_sva <= sigmoid_table_860_3_sva_dfm_1;
      sigmoid_table_859_0_sva <= sigmoid_table_859_0_sva_dfm_1;
      sigmoid_table_859_3_sva <= sigmoid_table_859_3_sva_dfm_1;
      sigmoid_table_858_0_sva <= sigmoid_table_858_0_sva_dfm_1;
      sigmoid_table_858_3_sva <= sigmoid_table_858_3_sva_dfm_1;
      sigmoid_table_857_0_sva <= sigmoid_table_857_0_sva_dfm_1;
      sigmoid_table_857_3_sva <= sigmoid_table_857_3_sva_dfm_1;
      sigmoid_table_856_0_sva <= sigmoid_table_856_0_sva_dfm_1;
      sigmoid_table_856_3_sva <= sigmoid_table_856_3_sva_dfm_1;
      sigmoid_table_855_0_sva <= sigmoid_table_855_0_sva_dfm_1;
      sigmoid_table_855_3_sva <= sigmoid_table_855_3_sva_dfm_1;
      sigmoid_table_854_0_sva <= sigmoid_table_854_0_sva_dfm_1;
      sigmoid_table_854_3_sva <= sigmoid_table_854_3_sva_dfm_1;
      sigmoid_table_853_0_sva <= sigmoid_table_853_0_sva_dfm_1;
      sigmoid_table_853_3_sva <= sigmoid_table_853_3_sva_dfm_1;
      sigmoid_table_852_3_sva <= sigmoid_table_852_3_sva_dfm_1;
      sigmoid_table_851_3_sva <= sigmoid_table_851_3_sva_dfm_1;
      sigmoid_table_850_3_sva <= sigmoid_table_850_3_sva_dfm_1;
      sigmoid_table_849_3_sva <= sigmoid_table_849_3_sva_dfm_1;
      sigmoid_table_848_3_sva <= sigmoid_table_848_3_sva_dfm_1;
      sigmoid_table_847_3_sva <= sigmoid_table_847_3_sva_dfm_1;
      sigmoid_table_846_3_sva <= sigmoid_table_846_3_sva_dfm_1;
      sigmoid_table_845_3_sva <= sigmoid_table_845_3_sva_dfm_1;
      sigmoid_table_844_3_sva <= sigmoid_table_844_3_sva_dfm_1;
      sigmoid_table_843_3_sva <= sigmoid_table_843_3_sva_dfm_1;
      sigmoid_table_842_3_sva <= sigmoid_table_842_3_sva_dfm_1;
      sigmoid_table_841_3_sva <= sigmoid_table_841_3_sva_dfm_1;
      sigmoid_table_840_3_sva <= sigmoid_table_840_3_sva_dfm_1;
      sigmoid_table_839_3_sva <= sigmoid_table_839_3_sva_dfm_1;
      sigmoid_table_838_3_sva <= sigmoid_table_838_3_sva_dfm_1;
      sigmoid_table_837_3_sva <= sigmoid_table_837_3_sva_dfm_1;
      sigmoid_table_836_3_sva <= sigmoid_table_836_3_sva_dfm_1;
      sigmoid_table_835_3_sva <= sigmoid_table_835_3_sva_dfm_1;
      sigmoid_table_834_3_sva <= sigmoid_table_834_3_sva_dfm_1;
      sigmoid_table_833_3_sva <= sigmoid_table_833_3_sva_dfm_1;
      sigmoid_table_832_3_sva <= sigmoid_table_832_3_sva_dfm_1;
      sigmoid_table_831_3_sva <= sigmoid_table_831_3_sva_dfm_1;
      sigmoid_table_830_3_sva <= sigmoid_table_830_3_sva_dfm_1;
      sigmoid_table_829_3_sva <= sigmoid_table_829_3_sva_dfm_1;
      sigmoid_table_828_3_sva <= sigmoid_table_828_3_sva_dfm_1;
      sigmoid_table_827_3_sva <= sigmoid_table_827_3_sva_dfm_1;
      sigmoid_table_826_3_sva <= sigmoid_table_826_3_sva_dfm_1;
      sigmoid_table_825_3_sva <= sigmoid_table_825_3_sva_dfm_1;
      sigmoid_table_824_3_sva <= sigmoid_table_824_3_sva_dfm_1;
      sigmoid_table_823_3_sva <= sigmoid_table_823_3_sva_dfm_1;
      sigmoid_table_822_3_sva <= sigmoid_table_822_3_sva_dfm_1;
      sigmoid_table_821_0_sva <= sigmoid_table_821_0_sva_dfm_1;
      sigmoid_table_821_4_sva <= sigmoid_table_821_4_sva_dfm_1;
      sigmoid_table_820_0_sva <= sigmoid_table_820_0_sva_dfm_1;
      sigmoid_table_820_4_sva <= sigmoid_table_820_4_sva_dfm_1;
      sigmoid_table_819_0_sva <= sigmoid_table_819_0_sva_dfm_1;
      sigmoid_table_819_4_sva <= sigmoid_table_819_4_sva_dfm_1;
      sigmoid_table_818_0_sva <= sigmoid_table_818_0_sva_dfm_1;
      sigmoid_table_818_4_sva <= sigmoid_table_818_4_sva_dfm_1;
      sigmoid_table_817_0_sva <= sigmoid_table_817_0_sva_dfm_1;
      sigmoid_table_817_4_sva <= sigmoid_table_817_4_sva_dfm_1;
      sigmoid_table_816_0_sva <= sigmoid_table_816_0_sva_dfm_1;
      sigmoid_table_816_4_sva <= sigmoid_table_816_4_sva_dfm_1;
      sigmoid_table_815_0_sva <= sigmoid_table_815_0_sva_dfm_1;
      sigmoid_table_815_4_sva <= sigmoid_table_815_4_sva_dfm_1;
      sigmoid_table_814_1_sva <= sigmoid_table_814_1_sva_dfm_1;
      sigmoid_table_814_4_sva <= sigmoid_table_814_4_sva_dfm_1;
      sigmoid_table_813_1_sva <= sigmoid_table_813_1_sva_dfm_1;
      sigmoid_table_813_4_sva <= sigmoid_table_813_4_sva_dfm_1;
      sigmoid_table_812_1_sva <= sigmoid_table_812_1_sva_dfm_1;
      sigmoid_table_812_4_sva <= sigmoid_table_812_4_sva_dfm_1;
      sigmoid_table_811_1_sva <= sigmoid_table_811_1_sva_dfm_1;
      sigmoid_table_811_4_sva <= sigmoid_table_811_4_sva_dfm_1;
      sigmoid_table_810_1_sva <= sigmoid_table_810_1_sva_dfm_1;
      sigmoid_table_810_4_sva <= sigmoid_table_810_4_sva_dfm_1;
      sigmoid_table_809_1_sva <= sigmoid_table_809_1_sva_dfm_1;
      sigmoid_table_809_4_sva <= sigmoid_table_809_4_sva_dfm_1;
      sigmoid_table_808_1_sva <= sigmoid_table_808_1_sva_dfm_1;
      sigmoid_table_808_4_sva <= sigmoid_table_808_4_sva_dfm_1;
      sigmoid_table_807_4_sva <= sigmoid_table_807_4_sva_dfm_1;
      sigmoid_table_806_4_sva <= sigmoid_table_806_4_sva_dfm_1;
      sigmoid_table_805_4_sva <= sigmoid_table_805_4_sva_dfm_1;
      sigmoid_table_804_4_sva <= sigmoid_table_804_4_sva_dfm_1;
      sigmoid_table_803_4_sva <= sigmoid_table_803_4_sva_dfm_1;
      sigmoid_table_802_4_sva <= sigmoid_table_802_4_sva_dfm_1;
      sigmoid_table_801_4_sva <= sigmoid_table_801_4_sva_dfm_1;
      sigmoid_table_800_4_sva <= sigmoid_table_800_4_sva_dfm_1;
      sigmoid_table_799_4_sva <= sigmoid_table_799_4_sva_dfm_1;
      sigmoid_table_798_4_sva <= sigmoid_table_798_4_sva_dfm_1;
      sigmoid_table_797_4_sva <= sigmoid_table_797_4_sva_dfm_1;
      sigmoid_table_796_4_sva <= sigmoid_table_796_4_sva_dfm_1;
      sigmoid_table_795_0_sva <= sigmoid_table_795_0_sva_dfm_1;
      sigmoid_table_795_4_sva <= sigmoid_table_795_4_sva_dfm_1;
      sigmoid_table_794_0_sva <= sigmoid_table_794_0_sva_dfm_1;
      sigmoid_table_794_4_sva <= sigmoid_table_794_4_sva_dfm_1;
      sigmoid_table_793_0_sva <= sigmoid_table_793_0_sva_dfm_1;
      sigmoid_table_793_4_sva <= sigmoid_table_793_4_sva_dfm_1;
      sigmoid_table_792_0_sva <= sigmoid_table_792_0_sva_dfm_1;
      sigmoid_table_792_4_sva <= sigmoid_table_792_4_sva_dfm_1;
      sigmoid_table_791_0_sva <= sigmoid_table_791_0_sva_dfm_1;
      sigmoid_table_791_4_sva <= sigmoid_table_791_4_sva_dfm_1;
      sigmoid_table_790_4_sva <= sigmoid_table_790_4_sva_dfm_1;
      sigmoid_table_789_4_sva <= sigmoid_table_789_4_sva_dfm_1;
      sigmoid_table_788_4_sva <= sigmoid_table_788_4_sva_dfm_1;
      sigmoid_table_787_4_sva <= sigmoid_table_787_4_sva_dfm_1;
      sigmoid_table_786_4_sva <= sigmoid_table_786_4_sva_dfm_1;
      sigmoid_table_785_4_sva <= sigmoid_table_785_4_sva_dfm_1;
      sigmoid_table_784_4_sva <= sigmoid_table_784_4_sva_dfm_1;
      sigmoid_table_783_4_sva <= sigmoid_table_783_4_sva_dfm_1;
      sigmoid_table_782_4_sva <= sigmoid_table_782_4_sva_dfm_1;
      sigmoid_table_781_4_sva <= sigmoid_table_781_4_sva_dfm_1;
      sigmoid_table_780_4_sva <= sigmoid_table_780_4_sva_dfm_1;
      sigmoid_table_779_4_sva <= sigmoid_table_779_4_sva_dfm_1;
      sigmoid_table_778_4_sva <= sigmoid_table_778_4_sva_dfm_1;
      sigmoid_table_777_0_sva <= sigmoid_table_777_0_sva_dfm_1;
      sigmoid_table_777_5_sva <= sigmoid_table_777_5_sva_dfm_1;
      sigmoid_table_776_0_sva <= sigmoid_table_776_0_sva_dfm_1;
      sigmoid_table_776_5_sva <= sigmoid_table_776_5_sva_dfm_1;
      sigmoid_table_775_0_sva <= sigmoid_table_775_0_sva_dfm_1;
      sigmoid_table_775_5_sva <= sigmoid_table_775_5_sva_dfm_1;
      sigmoid_table_774_0_sva <= sigmoid_table_774_0_sva_dfm_1;
      sigmoid_table_774_5_sva <= sigmoid_table_774_5_sva_dfm_1;
      sigmoid_table_773_1_sva <= sigmoid_table_773_1_sva_dfm_1;
      sigmoid_table_773_5_sva <= sigmoid_table_773_5_sva_dfm_1;
      sigmoid_table_772_1_sva <= sigmoid_table_772_1_sva_dfm_1;
      sigmoid_table_772_5_sva <= sigmoid_table_772_5_sva_dfm_1;
      sigmoid_table_771_1_sva <= sigmoid_table_771_1_sva_dfm_1;
      sigmoid_table_771_5_sva <= sigmoid_table_771_5_sva_dfm_1;
      sigmoid_table_770_1_sva <= sigmoid_table_770_1_sva_dfm_1;
      sigmoid_table_770_5_sva <= sigmoid_table_770_5_sva_dfm_1;
      sigmoid_table_769_2_sva <= sigmoid_table_769_2_sva_dfm_1;
      sigmoid_table_769_5_sva <= sigmoid_table_769_5_sva_dfm_1;
      sigmoid_table_768_2_sva <= sigmoid_table_768_2_sva_dfm_1;
      sigmoid_table_768_5_sva <= sigmoid_table_768_5_sva_dfm_1;
      sigmoid_table_767_2_sva <= sigmoid_table_767_2_sva_dfm_1;
      sigmoid_table_767_5_sva <= sigmoid_table_767_5_sva_dfm_1;
      sigmoid_table_766_2_sva <= sigmoid_table_766_2_sva_dfm_1;
      sigmoid_table_766_5_sva <= sigmoid_table_766_5_sva_dfm_1;
      sigmoid_table_765_2_sva <= sigmoid_table_765_2_sva_dfm_1;
      sigmoid_table_765_5_sva <= sigmoid_table_765_5_sva_dfm_1;
      sigmoid_table_764_2_sva <= sigmoid_table_764_2_sva_dfm_1;
      sigmoid_table_764_5_sva <= sigmoid_table_764_5_sva_dfm_1;
      sigmoid_table_763_2_sva <= sigmoid_table_763_2_sva_dfm_1;
      sigmoid_table_763_5_sva <= sigmoid_table_763_5_sva_dfm_1;
      sigmoid_table_762_0_sva <= sigmoid_table_762_0_sva_dfm_1;
      sigmoid_table_762_5_sva <= sigmoid_table_762_5_sva_dfm_1;
      sigmoid_table_761_0_sva <= sigmoid_table_761_0_sva_dfm_1;
      sigmoid_table_761_5_sva <= sigmoid_table_761_5_sva_dfm_1;
      sigmoid_table_760_0_sva <= sigmoid_table_760_0_sva_dfm_1;
      sigmoid_table_760_5_sva <= sigmoid_table_760_5_sva_dfm_1;
      sigmoid_table_759_5_sva <= sigmoid_table_759_5_sva_dfm_1;
      sigmoid_table_758_5_sva <= sigmoid_table_758_5_sva_dfm_1;
      sigmoid_table_757_5_sva <= sigmoid_table_757_5_sva_dfm_1;
      sigmoid_table_756_5_sva <= sigmoid_table_756_5_sva_dfm_1;
      sigmoid_table_755_5_sva <= sigmoid_table_755_5_sva_dfm_1;
      sigmoid_table_754_5_sva <= sigmoid_table_754_5_sva_dfm_1;
      sigmoid_table_753_5_sva <= sigmoid_table_753_5_sva_dfm_1;
      sigmoid_table_752_5_sva <= sigmoid_table_752_5_sva_dfm_1;
      sigmoid_table_751_5_sva <= sigmoid_table_751_5_sva_dfm_1;
      sigmoid_table_750_0_sva <= sigmoid_table_750_0_sva_dfm_1;
      sigmoid_table_750_5_sva <= sigmoid_table_750_5_sva_dfm_1;
      sigmoid_table_749_0_sva <= sigmoid_table_749_0_sva_dfm_1;
      sigmoid_table_749_5_sva <= sigmoid_table_749_5_sva_dfm_1;
      sigmoid_table_748_0_sva <= sigmoid_table_748_0_sva_dfm_1;
      sigmoid_table_748_5_sva <= sigmoid_table_748_5_sva_dfm_1;
      sigmoid_table_747_1_sva <= sigmoid_table_747_1_sva_dfm_1;
      sigmoid_table_747_5_sva <= sigmoid_table_747_5_sva_dfm_1;
      sigmoid_table_746_1_sva <= sigmoid_table_746_1_sva_dfm_1;
      sigmoid_table_746_5_sva <= sigmoid_table_746_5_sva_dfm_1;
      sigmoid_table_745_5_sva <= sigmoid_table_745_5_sva_dfm_1;
      sigmoid_table_744_5_sva <= sigmoid_table_744_5_sva_dfm_1;
      sigmoid_table_743_5_sva <= sigmoid_table_743_5_sva_dfm_1;
      sigmoid_table_742_5_sva <= sigmoid_table_742_5_sva_dfm_1;
      sigmoid_table_741_5_sva <= sigmoid_table_741_5_sva_dfm_1;
      sigmoid_table_740_0_sva <= sigmoid_table_740_0_sva_dfm_1;
      sigmoid_table_740_5_sva <= sigmoid_table_740_5_sva_dfm_1;
      sigmoid_table_739_0_sva <= sigmoid_table_739_0_sva_dfm_1;
      sigmoid_table_739_5_sva <= sigmoid_table_739_5_sva_dfm_1;
      sigmoid_table_738_5_sva <= sigmoid_table_738_5_sva_dfm_1;
      sigmoid_table_737_5_sva <= sigmoid_table_737_5_sva_dfm_1;
      sigmoid_table_736_5_sva <= sigmoid_table_736_5_sva_dfm_1;
      sigmoid_table_735_5_sva <= sigmoid_table_735_5_sva_dfm_1;
      sigmoid_table_734_5_sva <= sigmoid_table_734_5_sva_dfm_1;
      sigmoid_table_733_5_sva <= sigmoid_table_733_5_sva_dfm_1;
      sigmoid_table_732_5_sva <= sigmoid_table_732_5_sva_dfm_1;
      sigmoid_table_731_0_sva <= sigmoid_table_731_0_sva_dfm_1;
      sigmoid_table_731_6_sva <= sigmoid_table_731_6_sva_dfm_1;
      sigmoid_table_730_0_sva <= sigmoid_table_730_0_sva_dfm_1;
      sigmoid_table_730_6_sva <= sigmoid_table_730_6_sva_dfm_1;
      sigmoid_table_729_1_sva <= sigmoid_table_729_1_sva_dfm_1;
      sigmoid_table_729_6_sva <= sigmoid_table_729_6_sva_dfm_1;
      sigmoid_table_728_1_sva <= sigmoid_table_728_1_sva_dfm_1;
      sigmoid_table_728_6_sva <= sigmoid_table_728_6_sva_dfm_1;
      sigmoid_table_727_2_sva <= sigmoid_table_727_2_sva_dfm_1;
      sigmoid_table_727_6_sva <= sigmoid_table_727_6_sva_dfm_1;
      sigmoid_table_726_2_sva <= sigmoid_table_726_2_sva_dfm_1;
      sigmoid_table_726_6_sva <= sigmoid_table_726_6_sva_dfm_1;
      sigmoid_table_725_2_sva <= sigmoid_table_725_2_sva_dfm_1;
      sigmoid_table_725_6_sva <= sigmoid_table_725_6_sva_dfm_1;
      sigmoid_table_724_2_sva <= sigmoid_table_724_2_sva_dfm_1;
      sigmoid_table_724_6_sva <= sigmoid_table_724_6_sva_dfm_1;
      sigmoid_table_723_0_sva <= sigmoid_table_723_0_sva_dfm_1;
      sigmoid_table_723_3_sva <= sigmoid_table_723_3_sva_dfm_1;
      sigmoid_table_723_6_sva <= sigmoid_table_723_6_sva_dfm_1;
      sigmoid_table_722_3_sva <= sigmoid_table_722_3_sva_dfm_1;
      sigmoid_table_722_6_sva <= sigmoid_table_722_6_sva_dfm_1;
      sigmoid_table_721_3_sva <= sigmoid_table_721_3_sva_dfm_1;
      sigmoid_table_721_6_sva <= sigmoid_table_721_6_sva_dfm_1;
      sigmoid_table_720_3_sva <= sigmoid_table_720_3_sva_dfm_1;
      sigmoid_table_720_6_sva <= sigmoid_table_720_6_sva_dfm_1;
      sigmoid_table_719_3_sva <= sigmoid_table_719_3_sva_dfm_1;
      sigmoid_table_719_6_sva <= sigmoid_table_719_6_sva_dfm_1;
      sigmoid_table_718_3_sva <= sigmoid_table_718_3_sva_dfm_1;
      sigmoid_table_718_6_sva <= sigmoid_table_718_6_sva_dfm_1;
      sigmoid_table_717_3_sva <= sigmoid_table_717_3_sva_dfm_1;
      sigmoid_table_717_6_sva <= sigmoid_table_717_6_sva_dfm_1;
      sigmoid_table_716_0_sva <= sigmoid_table_716_0_sva_dfm_1;
      sigmoid_table_716_6_sva <= sigmoid_table_716_6_sva_dfm_1;
      sigmoid_table_715_1_sva <= sigmoid_table_715_1_sva_dfm_1;
      sigmoid_table_715_6_sva <= sigmoid_table_715_6_sva_dfm_1;
      sigmoid_table_714_1_sva <= sigmoid_table_714_1_sva_dfm_1;
      sigmoid_table_714_6_sva <= sigmoid_table_714_6_sva_dfm_1;
      sigmoid_table_713_6_sva <= sigmoid_table_713_6_sva_dfm_1;
      sigmoid_table_712_6_sva <= sigmoid_table_712_6_sva_dfm_1;
      sigmoid_table_711_6_sva <= sigmoid_table_711_6_sva_dfm_1;
      sigmoid_table_710_0_sva <= sigmoid_table_710_0_sva_dfm_1;
      sigmoid_table_710_6_sva <= sigmoid_table_710_6_sva_dfm_1;
      sigmoid_table_709_6_sva <= sigmoid_table_709_6_sva_dfm_1;
      sigmoid_table_708_6_sva <= sigmoid_table_708_6_sva_dfm_1;
      sigmoid_table_707_6_sva <= sigmoid_table_707_6_sva_dfm_1;
      sigmoid_table_706_6_sva <= sigmoid_table_706_6_sva_dfm_1;
      sigmoid_table_705_6_sva <= sigmoid_table_705_6_sva_dfm_1;
      sigmoid_table_704_0_sva <= sigmoid_table_704_0_sva_dfm_1;
      sigmoid_table_704_6_sva <= sigmoid_table_704_6_sva_dfm_1;
      sigmoid_table_703_1_sva <= sigmoid_table_703_1_sva_dfm_1;
      sigmoid_table_703_6_sva <= sigmoid_table_703_6_sva_dfm_1;
      sigmoid_table_702_2_sva <= sigmoid_table_702_2_sva_dfm_1;
      sigmoid_table_702_6_sva <= sigmoid_table_702_6_sva_dfm_1;
      sigmoid_table_701_2_sva <= sigmoid_table_701_2_sva_dfm_1;
      sigmoid_table_701_6_sva <= sigmoid_table_701_6_sva_dfm_1;
      sigmoid_table_700_2_sva <= sigmoid_table_700_2_sva_dfm_1;
      sigmoid_table_700_6_sva <= sigmoid_table_700_6_sva_dfm_1;
      sigmoid_table_699_0_sva <= sigmoid_table_699_0_sva_dfm_1;
      sigmoid_table_699_6_sva <= sigmoid_table_699_6_sva_dfm_1;
      sigmoid_table_698_6_sva <= sigmoid_table_698_6_sva_dfm_1;
      sigmoid_table_697_6_sva <= sigmoid_table_697_6_sva_dfm_1;
      sigmoid_table_696_6_sva <= sigmoid_table_696_6_sva_dfm_1;
      sigmoid_table_695_6_sva <= sigmoid_table_695_6_sva_dfm_1;
      sigmoid_table_694_0_sva <= sigmoid_table_694_0_sva_dfm_1;
      sigmoid_table_694_6_sva <= sigmoid_table_694_6_sva_dfm_1;
      sigmoid_table_693_1_sva <= sigmoid_table_693_1_sva_dfm_1;
      sigmoid_table_693_6_sva <= sigmoid_table_693_6_sva_dfm_1;
      sigmoid_table_692_6_sva <= sigmoid_table_692_6_sva_dfm_1;
      sigmoid_table_691_6_sva <= sigmoid_table_691_6_sva_dfm_1;
      sigmoid_table_690_6_sva <= sigmoid_table_690_6_sva_dfm_1;
      sigmoid_table_689_0_sva <= sigmoid_table_689_0_sva_dfm_1;
      sigmoid_table_689_6_sva <= sigmoid_table_689_6_sva_dfm_1;
      sigmoid_table_688_6_sva <= sigmoid_table_688_6_sva_dfm_1;
      sigmoid_table_687_6_sva <= sigmoid_table_687_6_sva_dfm_1;
      sigmoid_table_686_6_sva <= sigmoid_table_686_6_sva_dfm_1;
      sigmoid_table_685_0_sva <= sigmoid_table_685_0_sva_dfm_1;
      sigmoid_table_685_7_sva <= sigmoid_table_685_7_sva_dfm_1;
      sigmoid_table_684_1_sva <= sigmoid_table_684_1_sva_dfm_1;
      sigmoid_table_684_7_sva <= sigmoid_table_684_7_sva_dfm_1;
      sigmoid_table_683_2_sva <= sigmoid_table_683_2_sva_dfm_1;
      sigmoid_table_683_7_sva <= sigmoid_table_683_7_sva_dfm_1;
      sigmoid_table_682_2_sva <= sigmoid_table_682_2_sva_dfm_1;
      sigmoid_table_682_7_sva <= sigmoid_table_682_7_sva_dfm_1;
      sigmoid_table_681_0_sva <= sigmoid_table_681_0_sva_dfm_1;
      sigmoid_table_681_3_sva <= sigmoid_table_681_3_sva_dfm_1;
      sigmoid_table_681_7_sva <= sigmoid_table_681_7_sva_dfm_1;
      sigmoid_table_680_3_sva <= sigmoid_table_680_3_sva_dfm_1;
      sigmoid_table_680_7_sva <= sigmoid_table_680_7_sva_dfm_1;
      sigmoid_table_679_3_sva <= sigmoid_table_679_3_sva_dfm_1;
      sigmoid_table_679_7_sva <= sigmoid_table_679_7_sva_dfm_1;
      sigmoid_table_678_3_sva <= sigmoid_table_678_3_sva_dfm_1;
      sigmoid_table_678_7_sva <= sigmoid_table_678_7_sva_dfm_1;
      sigmoid_table_677_0_sva <= sigmoid_table_677_0_sva_dfm_1;
      sigmoid_table_677_4_sva <= sigmoid_table_677_4_sva_dfm_1;
      sigmoid_table_677_7_sva <= sigmoid_table_677_7_sva_dfm_1;
      sigmoid_table_676_1_sva <= sigmoid_table_676_1_sva_dfm_1;
      sigmoid_table_676_4_sva <= sigmoid_table_676_4_sva_dfm_1;
      sigmoid_table_676_7_sva <= sigmoid_table_676_7_sva_dfm_1;
      sigmoid_table_675_4_sva <= sigmoid_table_675_4_sva_dfm_1;
      sigmoid_table_675_7_sva <= sigmoid_table_675_7_sva_dfm_1;
      sigmoid_table_674_4_sva <= sigmoid_table_674_4_sva_dfm_1;
      sigmoid_table_674_7_sva <= sigmoid_table_674_7_sva_dfm_1;
      sigmoid_table_673_0_sva <= sigmoid_table_673_0_sva_dfm_1;
      sigmoid_table_673_4_sva <= sigmoid_table_673_4_sva_dfm_1;
      sigmoid_table_673_7_sva <= sigmoid_table_673_7_sva_dfm_1;
      sigmoid_table_672_4_sva <= sigmoid_table_672_4_sva_dfm_1;
      sigmoid_table_672_7_sva <= sigmoid_table_672_7_sva_dfm_1;
      sigmoid_table_671_4_sva <= sigmoid_table_671_4_sva_dfm_1;
      sigmoid_table_671_7_sva <= sigmoid_table_671_7_sva_dfm_1;
      sigmoid_table_670_4_sva <= sigmoid_table_670_4_sva_dfm_1;
      sigmoid_table_670_7_sva <= sigmoid_table_670_7_sva_dfm_1;
      sigmoid_table_669_1_sva <= sigmoid_table_669_1_sva_dfm_1;
      sigmoid_table_669_7_sva <= sigmoid_table_669_7_sva_dfm_1;
      sigmoid_table_668_2_sva <= sigmoid_table_668_2_sva_dfm_1;
      sigmoid_table_668_7_sva <= sigmoid_table_668_7_sva_dfm_1;
      sigmoid_table_667_2_sva <= sigmoid_table_667_2_sva_dfm_1;
      sigmoid_table_667_7_sva <= sigmoid_table_667_7_sva_dfm_1;
      sigmoid_table_666_0_sva <= sigmoid_table_666_0_sva_dfm_1;
      sigmoid_table_666_7_sva <= sigmoid_table_666_7_sva_dfm_1;
      sigmoid_table_665_7_sva <= sigmoid_table_665_7_sva_dfm_1;
      sigmoid_table_664_7_sva <= sigmoid_table_664_7_sva_dfm_1;
      sigmoid_table_663_0_sva <= sigmoid_table_663_0_sva_dfm_1;
      sigmoid_table_663_7_sva <= sigmoid_table_663_7_sva_dfm_1;
      sigmoid_table_662_1_sva <= sigmoid_table_662_1_sva_dfm_1;
      sigmoid_table_662_7_sva <= sigmoid_table_662_7_sva_dfm_1;
      sigmoid_table_661_7_sva <= sigmoid_table_661_7_sva_dfm_1;
      sigmoid_table_660_0_sva <= sigmoid_table_660_0_sva_dfm_1;
      sigmoid_table_660_7_sva <= sigmoid_table_660_7_sva_dfm_1;
      sigmoid_table_659_7_sva <= sigmoid_table_659_7_sva_dfm_1;
      sigmoid_table_658_7_sva <= sigmoid_table_658_7_sva_dfm_1;
      sigmoid_table_657_0_sva <= sigmoid_table_657_0_sva_dfm_1;
      sigmoid_table_657_7_sva <= sigmoid_table_657_7_sva_dfm_1;
      sigmoid_table_656_1_sva <= sigmoid_table_656_1_sva_dfm_1;
      sigmoid_table_656_7_sva <= sigmoid_table_656_7_sva_dfm_1;
      sigmoid_table_655_2_sva <= sigmoid_table_655_2_sva_dfm_1;
      sigmoid_table_655_7_sva <= sigmoid_table_655_7_sva_dfm_1;
      sigmoid_table_654_0_sva <= sigmoid_table_654_0_sva_dfm_1;
      sigmoid_table_654_3_sva <= sigmoid_table_654_3_sva_dfm_1;
      sigmoid_table_654_7_sva <= sigmoid_table_654_7_sva_dfm_1;
      sigmoid_table_653_3_sva <= sigmoid_table_653_3_sva_dfm_1;
      sigmoid_table_653_7_sva <= sigmoid_table_653_7_sva_dfm_1;
      sigmoid_table_652_3_sva <= sigmoid_table_652_3_sva_dfm_1;
      sigmoid_table_652_7_sva <= sigmoid_table_652_7_sva_dfm_1;
      sigmoid_table_651_0_sva <= sigmoid_table_651_0_sva_dfm_1;
      sigmoid_table_651_7_sva <= sigmoid_table_651_7_sva_dfm_1;
      sigmoid_table_650_7_sva <= sigmoid_table_650_7_sva_dfm_1;
      sigmoid_table_649_7_sva <= sigmoid_table_649_7_sva_dfm_1;
      sigmoid_table_648_7_sva <= sigmoid_table_648_7_sva_dfm_1;
      sigmoid_table_647_7_sva <= sigmoid_table_647_7_sva_dfm_1;
      sigmoid_table_646_0_sva <= sigmoid_table_646_0_sva_dfm_1;
      sigmoid_table_646_7_sva <= sigmoid_table_646_7_sva_dfm_1;
      sigmoid_table_645_1_sva <= sigmoid_table_645_1_sva_dfm_1;
      sigmoid_table_645_7_sva <= sigmoid_table_645_7_sva_dfm_1;
      sigmoid_table_644_2_sva <= sigmoid_table_644_2_sva_dfm_1;
      sigmoid_table_644_7_sva <= sigmoid_table_644_7_sva_dfm_1;
      sigmoid_table_643_7_sva <= sigmoid_table_643_7_sva_dfm_1;
      sigmoid_table_642_7_sva <= sigmoid_table_642_7_sva_dfm_1;
      sigmoid_table_641_0_sva <= sigmoid_table_641_0_sva_dfm_1;
      sigmoid_table_641_7_sva <= sigmoid_table_641_7_sva_dfm_1;
      sigmoid_table_640_7_sva <= sigmoid_table_640_7_sva_dfm_1;
      sigmoid_table_639_7_sva <= sigmoid_table_639_7_sva_dfm_1;
      sigmoid_table_638_7_sva <= sigmoid_table_638_7_sva_dfm_1;
      sigmoid_table_637_7_sva <= sigmoid_table_637_7_sva_dfm_1;
      sigmoid_table_636_0_sva <= sigmoid_table_636_0_sva_dfm_1;
      sigmoid_table_636_8_sva <= sigmoid_table_636_8_sva_dfm_1;
      sigmoid_table_635_2_sva <= sigmoid_table_635_2_sva_dfm_1;
      sigmoid_table_635_8_sva <= sigmoid_table_635_8_sva_dfm_1;
      sigmoid_table_634_0_sva <= sigmoid_table_634_0_sva_dfm_1;
      sigmoid_table_634_3_sva <= sigmoid_table_634_3_sva_dfm_1;
      sigmoid_table_634_8_sva <= sigmoid_table_634_8_sva_dfm_1;
      sigmoid_table_633_3_sva <= sigmoid_table_633_3_sva_dfm_1;
      sigmoid_table_633_8_sva <= sigmoid_table_633_8_sva_dfm_1;
      sigmoid_table_632_0_sva <= sigmoid_table_632_0_sva_dfm_1;
      sigmoid_table_632_4_sva <= sigmoid_table_632_4_sva_dfm_1;
      sigmoid_table_632_8_sva <= sigmoid_table_632_8_sva_dfm_1;
      sigmoid_table_631_4_sva <= sigmoid_table_631_4_sva_dfm_1;
      sigmoid_table_631_8_sva <= sigmoid_table_631_8_sva_dfm_1;
      sigmoid_table_630_4_sva <= sigmoid_table_630_4_sva_dfm_1;
      sigmoid_table_630_8_sva <= sigmoid_table_630_8_sva_dfm_1;
      sigmoid_table_629_4_sva <= sigmoid_table_629_4_sva_dfm_1;
      sigmoid_table_629_8_sva <= sigmoid_table_629_8_sva_dfm_1;
      sigmoid_table_628_4_sva <= sigmoid_table_628_4_sva_dfm_1;
      sigmoid_table_628_8_sva <= sigmoid_table_628_8_sva_dfm_1;
      sigmoid_table_627_1_sva <= sigmoid_table_627_1_sva_dfm_1;
      sigmoid_table_627_5_sva <= sigmoid_table_627_5_sva_dfm_1;
      sigmoid_table_627_8_sva <= sigmoid_table_627_8_sva_dfm_1;
      sigmoid_table_626_2_sva <= sigmoid_table_626_2_sva_dfm_1;
      sigmoid_table_626_5_sva <= sigmoid_table_626_5_sva_dfm_1;
      sigmoid_table_626_8_sva <= sigmoid_table_626_8_sva_dfm_1;
      sigmoid_table_625_5_sva <= sigmoid_table_625_5_sva_dfm_1;
      sigmoid_table_625_8_sva <= sigmoid_table_625_8_sva_dfm_1;
      sigmoid_table_624_5_sva <= sigmoid_table_624_5_sva_dfm_1;
      sigmoid_table_624_8_sva <= sigmoid_table_624_8_sva_dfm_1;
      sigmoid_table_623_1_sva <= sigmoid_table_623_1_sva_dfm_1;
      sigmoid_table_623_5_sva <= sigmoid_table_623_5_sva_dfm_1;
      sigmoid_table_623_8_sva <= sigmoid_table_623_8_sva_dfm_1;
      sigmoid_table_622_5_sva <= sigmoid_table_622_5_sva_dfm_1;
      sigmoid_table_622_8_sva <= sigmoid_table_622_8_sva_dfm_1;
      sigmoid_table_621_5_sva <= sigmoid_table_621_5_sva_dfm_1;
      sigmoid_table_621_8_sva <= sigmoid_table_621_8_sva_dfm_1;
      sigmoid_table_620_5_sva <= sigmoid_table_620_5_sva_dfm_1;
      sigmoid_table_620_8_sva <= sigmoid_table_620_8_sva_dfm_1;
      sigmoid_table_619_1_sva <= sigmoid_table_619_1_sva_dfm_1;
      sigmoid_table_619_8_sva <= sigmoid_table_619_8_sva_dfm_1;
      sigmoid_table_618_0_sva <= sigmoid_table_618_0_sva_dfm_1;
      sigmoid_table_618_3_sva <= sigmoid_table_618_3_sva_dfm_1;
      sigmoid_table_618_8_sva <= sigmoid_table_618_8_sva_dfm_1;
      sigmoid_table_617_3_sva <= sigmoid_table_617_3_sva_dfm_1;
      sigmoid_table_617_8_sva <= sigmoid_table_617_8_sva_dfm_1;
      sigmoid_table_616_0_sva <= sigmoid_table_616_0_sva_dfm_1;
      sigmoid_table_616_8_sva <= sigmoid_table_616_8_sva_dfm_1;
      sigmoid_table_615_8_sva <= sigmoid_table_615_8_sva_dfm_1;
      sigmoid_table_614_0_sva <= sigmoid_table_614_0_sva_dfm_1;
      sigmoid_table_614_8_sva <= sigmoid_table_614_8_sva_dfm_1;
      sigmoid_table_613_8_sva <= sigmoid_table_613_8_sva_dfm_1;
      sigmoid_table_612_1_sva <= sigmoid_table_612_1_sva_dfm_1;
      sigmoid_table_612_8_sva <= sigmoid_table_612_8_sva_dfm_1;
      sigmoid_table_611_2_sva <= sigmoid_table_611_2_sva_dfm_1;
      sigmoid_table_611_8_sva <= sigmoid_table_611_8_sva_dfm_1;
      sigmoid_table_610_8_sva <= sigmoid_table_610_8_sva_dfm_1;
      sigmoid_table_609_0_sva <= sigmoid_table_609_0_sva_dfm_1;
      sigmoid_table_609_8_sva <= sigmoid_table_609_8_sva_dfm_1;
      sigmoid_table_608_8_sva <= sigmoid_table_608_8_sva_dfm_1;
      sigmoid_table_607_8_sva <= sigmoid_table_607_8_sva_dfm_1;
      sigmoid_table_606_8_sva <= sigmoid_table_606_8_sva_dfm_1;
      sigmoid_table_605_2_sva <= sigmoid_table_605_2_sva_dfm_1;
      sigmoid_table_605_8_sva <= sigmoid_table_605_8_sva_dfm_1;
      sigmoid_table_604_0_sva <= sigmoid_table_604_0_sva_dfm_1;
      sigmoid_table_604_3_sva <= sigmoid_table_604_3_sva_dfm_1;
      sigmoid_table_604_8_sva <= sigmoid_table_604_8_sva_dfm_1;
      sigmoid_table_603_3_sva <= sigmoid_table_603_3_sva_dfm_1;
      sigmoid_table_603_8_sva <= sigmoid_table_603_8_sva_dfm_1;
      sigmoid_table_602_1_sva <= sigmoid_table_602_1_sva_dfm_1;
      sigmoid_table_602_4_sva <= sigmoid_table_602_4_sva_dfm_1;
      sigmoid_table_602_8_sva <= sigmoid_table_602_8_sva_dfm_1;
      sigmoid_table_601_0_sva <= sigmoid_table_601_0_sva_dfm_1;
      sigmoid_table_601_4_sva <= sigmoid_table_601_4_sva_dfm_1;
      sigmoid_table_601_8_sva <= sigmoid_table_601_8_sva_dfm_1;
      sigmoid_table_600_4_sva <= sigmoid_table_600_4_sva_dfm_1;
      sigmoid_table_600_8_sva <= sigmoid_table_600_8_sva_dfm_1;
      sigmoid_table_599_1_sva <= sigmoid_table_599_1_sva_dfm_1;
      sigmoid_table_599_8_sva <= sigmoid_table_599_8_sva_dfm_1;
      sigmoid_table_598_2_sva <= sigmoid_table_598_2_sva_dfm_1;
      sigmoid_table_598_8_sva <= sigmoid_table_598_8_sva_dfm_1;
      sigmoid_table_597_8_sva <= sigmoid_table_597_8_sva_dfm_1;
      sigmoid_table_596_1_sva <= sigmoid_table_596_1_sva_dfm_1;
      sigmoid_table_596_8_sva <= sigmoid_table_596_8_sva_dfm_1;
      sigmoid_table_595_8_sva <= sigmoid_table_595_8_sva_dfm_1;
      sigmoid_table_594_8_sva <= sigmoid_table_594_8_sva_dfm_1;
      sigmoid_table_593_1_sva <= sigmoid_table_593_1_sva_dfm_1;
      sigmoid_table_593_8_sva <= sigmoid_table_593_8_sva_dfm_1;
      sigmoid_table_592_0_sva <= sigmoid_table_592_0_sva_dfm_1;
      sigmoid_table_592_3_sva <= sigmoid_table_592_3_sva_dfm_1;
      sigmoid_table_592_8_sva <= sigmoid_table_592_8_sva_dfm_1;
      sigmoid_table_591_3_sva <= sigmoid_table_591_3_sva_dfm_1;
      sigmoid_table_591_8_sva <= sigmoid_table_591_8_sva_dfm_1;
      sigmoid_table_590_1_sva <= sigmoid_table_590_1_sva_dfm_1;
      sigmoid_table_590_8_sva <= sigmoid_table_590_8_sva_dfm_1;
      sigmoid_table_589_0_sva <= sigmoid_table_589_0_sva_dfm_1;
      sigmoid_table_589_8_sva <= sigmoid_table_589_8_sva_dfm_1;
      sigmoid_table_588_8_sva <= sigmoid_table_588_8_sva_dfm_1;
      sigmoid_table_587_2_sva <= sigmoid_table_587_2_sva_dfm_1;
      sigmoid_table_587_8_sva <= sigmoid_table_587_8_sva_dfm_1;
      sigmoid_table_586_8_sva <= sigmoid_table_586_8_sva_dfm_1;
      sigmoid_table_585_0_sva <= sigmoid_table_585_0_sva_dfm_1;
      sigmoid_table_585_8_sva <= sigmoid_table_585_8_sva_dfm_1;
      sigmoid_table_584_8_sva <= sigmoid_table_584_8_sva_dfm_1;
      sigmoid_table_583_8_sva <= sigmoid_table_583_8_sva_dfm_1;
      sigmoid_table_582_0_sva <= sigmoid_table_582_0_sva_dfm_1;
      sigmoid_table_581_2_sva <= sigmoid_table_581_2_sva_dfm_1;
      sigmoid_table_580_3_sva <= sigmoid_table_580_3_sva_dfm_1;
      sigmoid_table_579_4_sva <= sigmoid_table_579_4_sva_dfm_1;
      sigmoid_table_578_4_sva <= sigmoid_table_578_4_sva_dfm_1;
      sigmoid_table_577_0_sva <= sigmoid_table_577_0_sva_dfm_1;
      sigmoid_table_577_5_sva <= sigmoid_table_577_5_sva_dfm_1;
      sigmoid_table_576_2_sva <= sigmoid_table_576_2_sva_dfm_1;
      sigmoid_table_576_5_sva <= sigmoid_table_576_5_sva_dfm_1;
      sigmoid_table_575_5_sva <= sigmoid_table_575_5_sva_dfm_1;
      sigmoid_table_574_1_sva <= sigmoid_table_574_1_sva_dfm_1;
      sigmoid_table_574_5_sva <= sigmoid_table_574_5_sva_dfm_1;
      sigmoid_table_573_0_sva <= sigmoid_table_573_0_sva_dfm_1;
      sigmoid_table_573_5_sva <= sigmoid_table_573_5_sva_dfm_1;
      sigmoid_table_572_0_sva <= sigmoid_table_572_0_sva_dfm_1;
      sigmoid_table_572_6_sva <= sigmoid_table_572_6_sva_dfm_1;
      sigmoid_table_571_2_sva <= sigmoid_table_571_2_sva_dfm_1;
      sigmoid_table_571_6_sva <= sigmoid_table_571_6_sva_dfm_1;
      sigmoid_table_570_3_sva <= sigmoid_table_570_3_sva_dfm_1;
      sigmoid_table_570_6_sva <= sigmoid_table_570_6_sva_dfm_1;
      sigmoid_table_569_1_sva <= sigmoid_table_569_1_sva_dfm_1;
      sigmoid_table_569_6_sva <= sigmoid_table_569_6_sva_dfm_1;
      sigmoid_table_568_6_sva <= sigmoid_table_568_6_sva_dfm_1;
      sigmoid_table_567_0_sva <= sigmoid_table_567_0_sva_dfm_1;
      sigmoid_table_567_6_sva <= sigmoid_table_567_6_sva_dfm_1;
      sigmoid_table_566_2_sva <= sigmoid_table_566_2_sva_dfm_1;
      sigmoid_table_566_6_sva <= sigmoid_table_566_6_sva_dfm_1;
      sigmoid_table_565_6_sva <= sigmoid_table_565_6_sva_dfm_1;
      sigmoid_table_564_6_sva <= sigmoid_table_564_6_sva_dfm_1;
      sigmoid_table_563_6_sva <= sigmoid_table_563_6_sva_dfm_1;
      sigmoid_table_562_1_sva <= sigmoid_table_562_1_sva_dfm_1;
      sigmoid_table_561_3_sva <= sigmoid_table_561_3_sva_dfm_1;
      sigmoid_table_560_0_sva <= sigmoid_table_560_0_sva_dfm_1;
      sigmoid_table_560_4_sva <= sigmoid_table_560_4_sva_dfm_1;
      sigmoid_table_559_0_sva <= sigmoid_table_559_0_sva_dfm_1;
      sigmoid_table_559_4_sva <= sigmoid_table_559_4_sva_dfm_1;
      sigmoid_table_558_4_sva <= sigmoid_table_558_4_sva_dfm_1;
      sigmoid_table_557_2_sva <= sigmoid_table_557_2_sva_dfm_1;
      sigmoid_table_553_1_sva <= sigmoid_table_553_1_sva_dfm_1;
      sigmoid_table_552_3_sva <= sigmoid_table_552_3_sva_dfm_1;
      sigmoid_table_551_0_sva <= sigmoid_table_551_0_sva_dfm_1;
      sigmoid_table_550_0_sva <= sigmoid_table_550_0_sva_dfm_1;
      sigmoid_table_548_2_sva <= sigmoid_table_548_2_sva_dfm_1;
      sigmoid_table_544_2_sva <= sigmoid_table_544_2_sva_dfm_1;
      sigmoid_table_543_3_sva <= sigmoid_table_543_3_sva_dfm_1;
      sigmoid_table_542_4_sva <= sigmoid_table_542_4_sva_dfm_1;
      sigmoid_table_541_4_sva <= sigmoid_table_541_4_sva_dfm_1;
      sigmoid_table_540_1_sva <= sigmoid_table_540_1_sva_dfm_1;
      sigmoid_table_540_5_sva <= sigmoid_table_540_5_sva_dfm_1;
      sigmoid_table_539_5_sva <= sigmoid_table_539_5_sva_dfm_1;
      sigmoid_table_538_1_sva <= sigmoid_table_538_1_sva_dfm_1;
      sigmoid_table_538_5_sva <= sigmoid_table_538_5_sva_dfm_1;
      sigmoid_table_537_5_sva <= sigmoid_table_537_5_sva_dfm_1;
      sigmoid_table_536_1_sva <= sigmoid_table_536_1_sva_dfm_1;
      sigmoid_table_535_0_sva <= sigmoid_table_535_0_sva_dfm_1;
      sigmoid_table_535_3_sva <= sigmoid_table_535_3_sva_dfm_1;
      sigmoid_table_534_0_sva <= sigmoid_table_534_0_sva_dfm_1;
      sigmoid_table_533_0_sva <= sigmoid_table_533_0_sva_dfm_1;
      sigmoid_table_532_0_sva <= sigmoid_table_532_0_sva_dfm_1;
      sigmoid_table_531_0_sva <= sigmoid_table_531_0_sva_dfm_1;
      sigmoid_table_530_0_sva <= sigmoid_table_530_0_sva_dfm_1;
      sigmoid_table_529_0_sva <= sigmoid_table_529_0_sva_dfm_1;
      sigmoid_table_528_0_sva <= sigmoid_table_528_0_sva_dfm_1;
      sigmoid_table_527_0_sva <= sigmoid_table_527_0_sva_dfm_1;
      sigmoid_table_527_3_sva <= sigmoid_table_527_3_sva_dfm_1;
      sigmoid_table_526_0_sva <= sigmoid_table_526_0_sva_dfm_1;
      sigmoid_table_526_4_sva <= sigmoid_table_526_4_sva_dfm_1;
      sigmoid_table_525_0_sva <= sigmoid_table_525_0_sva_dfm_1;
      sigmoid_table_525_4_sva <= sigmoid_table_525_4_sva_dfm_1;
      sigmoid_table_524_0_sva <= sigmoid_table_524_0_sva_dfm_1;
      sigmoid_table_523_0_sva <= sigmoid_table_523_0_sva_dfm_1;
      sigmoid_table_522_0_sva <= sigmoid_table_522_0_sva_dfm_1;
      sigmoid_table_521_0_sva <= sigmoid_table_521_0_sva_dfm_1;
      sigmoid_table_520_0_sva <= sigmoid_table_520_0_sva_dfm_1;
      sigmoid_table_519_0_sva <= sigmoid_table_519_0_sva_dfm_1;
      sigmoid_table_519_3_sva <= sigmoid_table_519_3_sva_dfm_1;
      sigmoid_table_518_0_sva <= sigmoid_table_518_0_sva_dfm_1;
      sigmoid_table_517_0_sva <= sigmoid_table_517_0_sva_dfm_1;
      sigmoid_table_516_0_sva <= sigmoid_table_516_0_sva_dfm_1;
      sigmoid_table_515_2_sva <= sigmoid_table_515_2_sva_dfm_1;
      sigmoid_table_511_2_sva <= sigmoid_table_511_2_sva_dfm_1;
      sigmoid_table_510_3_sva <= sigmoid_table_510_3_sva_dfm_1;
      sigmoid_table_509_4_sva <= sigmoid_table_509_4_sva_dfm_1;
      sigmoid_table_508_4_sva <= sigmoid_table_508_4_sva_dfm_1;
      sigmoid_table_507_2_sva <= sigmoid_table_507_2_sva_dfm_1;
      sigmoid_table_507_5_sva <= sigmoid_table_507_5_sva_dfm_1;
      sigmoid_table_506_5_sva <= sigmoid_table_506_5_sva_dfm_1;
      sigmoid_table_505_5_sva <= sigmoid_table_505_5_sva_dfm_1;
      sigmoid_table_504_5_sva <= sigmoid_table_504_5_sva_dfm_1;
      sigmoid_table_503_2_sva <= sigmoid_table_503_2_sva_dfm_1;
      sigmoid_table_503_6_sva <= sigmoid_table_503_6_sva_dfm_1;
      sigmoid_table_502_3_sva <= sigmoid_table_502_3_sva_dfm_1;
      sigmoid_table_502_6_sva <= sigmoid_table_502_6_sva_dfm_1;
      sigmoid_table_501_6_sva <= sigmoid_table_501_6_sva_dfm_1;
      sigmoid_table_500_6_sva <= sigmoid_table_500_6_sva_dfm_1;
      sigmoid_table_499_2_sva <= sigmoid_table_499_2_sva_dfm_1;
      sigmoid_table_499_6_sva <= sigmoid_table_499_6_sva_dfm_1;
      sigmoid_table_498_6_sva <= sigmoid_table_498_6_sva_dfm_1;
      sigmoid_table_497_6_sva <= sigmoid_table_497_6_sva_dfm_1;
      sigmoid_table_496_6_sva <= sigmoid_table_496_6_sva_dfm_1;
      sigmoid_table_495_2_sva <= sigmoid_table_495_2_sva_dfm_1;
      sigmoid_table_495_7_sva <= sigmoid_table_495_7_sva_dfm_1;
      sigmoid_table_494_3_sva <= sigmoid_table_494_3_sva_dfm_1;
      sigmoid_table_494_7_sva <= sigmoid_table_494_7_sva_dfm_1;
      sigmoid_table_493_4_sva <= sigmoid_table_493_4_sva_dfm_1;
      sigmoid_table_493_7_sva <= sigmoid_table_493_7_sva_dfm_1;
      sigmoid_table_492_4_sva <= sigmoid_table_492_4_sva_dfm_1;
      sigmoid_table_492_7_sva <= sigmoid_table_492_7_sva_dfm_1;
      sigmoid_table_491_2_sva <= sigmoid_table_491_2_sva_dfm_1;
      sigmoid_table_491_7_sva <= sigmoid_table_491_7_sva_dfm_1;
      sigmoid_table_490_7_sva <= sigmoid_table_490_7_sva_dfm_1;
      sigmoid_table_489_7_sva <= sigmoid_table_489_7_sva_dfm_1;
      sigmoid_table_488_7_sva <= sigmoid_table_488_7_sva_dfm_1;
      sigmoid_table_487_2_sva <= sigmoid_table_487_2_sva_dfm_1;
      sigmoid_table_487_7_sva <= sigmoid_table_487_7_sva_dfm_1;
      sigmoid_table_486_3_sva <= sigmoid_table_486_3_sva_dfm_1;
      sigmoid_table_486_7_sva <= sigmoid_table_486_7_sva_dfm_1;
      sigmoid_table_485_7_sva <= sigmoid_table_485_7_sva_dfm_1;
      sigmoid_table_484_7_sva <= sigmoid_table_484_7_sva_dfm_1;
      sigmoid_table_483_2_sva <= sigmoid_table_483_2_sva_dfm_1;
      sigmoid_table_483_7_sva <= sigmoid_table_483_7_sva_dfm_1;
      sigmoid_table_482_7_sva <= sigmoid_table_482_7_sva_dfm_1;
      sigmoid_table_481_1_sva <= sigmoid_table_481_1_sva_dfm_1;
      sigmoid_table_481_7_sva <= sigmoid_table_481_7_sva_dfm_1;
      sigmoid_table_480_7_sva <= sigmoid_table_480_7_sva_dfm_1;
      sigmoid_table_479_1_sva <= sigmoid_table_479_1_sva_dfm_1;
      sigmoid_table_478_0_sva <= sigmoid_table_478_0_sva_dfm_1;
      sigmoid_table_478_3_sva <= sigmoid_table_478_3_sva_dfm_1;
      sigmoid_table_477_0_sva <= sigmoid_table_477_0_sva_dfm_1;
      sigmoid_table_477_4_sva <= sigmoid_table_477_4_sva_dfm_1;
      sigmoid_table_476_0_sva <= sigmoid_table_476_0_sva_dfm_1;
      sigmoid_table_476_4_sva <= sigmoid_table_476_4_sva_dfm_1;
      sigmoid_table_475_0_sva <= sigmoid_table_475_0_sva_dfm_1;
      sigmoid_table_475_5_sva <= sigmoid_table_475_5_sva_dfm_1;
      sigmoid_table_474_2_sva <= sigmoid_table_474_2_sva_dfm_1;
      sigmoid_table_474_5_sva <= sigmoid_table_474_5_sva_dfm_1;
      sigmoid_table_473_5_sva <= sigmoid_table_473_5_sva_dfm_1;
      sigmoid_table_472_5_sva <= sigmoid_table_472_5_sva_dfm_1;
      sigmoid_table_471_5_sva <= sigmoid_table_471_5_sva_dfm_1;
      sigmoid_table_470_2_sva <= sigmoid_table_470_2_sva_dfm_1;
      sigmoid_table_469_3_sva <= sigmoid_table_469_3_sva_dfm_1;
      sigmoid_table_468_1_sva <= sigmoid_table_468_1_sva_dfm_1;
      sigmoid_table_467_0_sva <= sigmoid_table_467_0_sva_dfm_1;
      sigmoid_table_466_0_sva <= sigmoid_table_466_0_sva_dfm_1;
      sigmoid_table_465_2_sva <= sigmoid_table_465_2_sva_dfm_1;
      sigmoid_table_461_1_sva <= sigmoid_table_461_1_sva_dfm_1;
      sigmoid_table_460_3_sva <= sigmoid_table_460_3_sva_dfm_1;
      sigmoid_table_459_0_sva <= sigmoid_table_459_0_sva_dfm_1;
      sigmoid_table_459_4_sva <= sigmoid_table_459_4_sva_dfm_1;
      sigmoid_table_458_0_sva <= sigmoid_table_458_0_sva_dfm_1;
      sigmoid_table_458_4_sva <= sigmoid_table_458_4_sva_dfm_1;
      sigmoid_table_457_4_sva <= sigmoid_table_457_4_sva_dfm_1;
      sigmoid_table_456_2_sva <= sigmoid_table_456_2_sva_dfm_1;
      sigmoid_table_454_1_sva <= sigmoid_table_454_1_sva_dfm_1;
      sigmoid_table_453_0_sva <= sigmoid_table_453_0_sva_dfm_1;
      sigmoid_table_451_2_sva <= sigmoid_table_451_2_sva_dfm_1;
      sigmoid_table_450_3_sva <= sigmoid_table_450_3_sva_dfm_1;
      sigmoid_table_449_1_sva <= sigmoid_table_449_1_sva_dfm_1;
      sigmoid_table_448_0_sva <= sigmoid_table_448_0_sva_dfm_1;
      sigmoid_table_446_2_sva <= sigmoid_table_446_2_sva_dfm_1;
      sigmoid_table_444_1_sva <= sigmoid_table_444_1_sva_dfm_1;
      sigmoid_table_443_0_sva <= sigmoid_table_443_0_sva_dfm_1;
      sigmoid_table_441_2_sva <= sigmoid_table_441_2_sva_dfm_1;
      sigmoid_table_440_3_sva <= sigmoid_table_440_3_sva_dfm_1;
      sigmoid_table_439_3_sva <= sigmoid_table_439_3_sva_dfm_1;
      sigmoid_table_438_4_sva <= sigmoid_table_438_4_sva_dfm_1;
      sigmoid_table_437_4_sva <= sigmoid_table_437_4_sva_dfm_1;
      sigmoid_table_436_0_sva <= sigmoid_table_436_0_sva_dfm_1;
      sigmoid_table_436_5_sva <= sigmoid_table_436_5_sva_dfm_1;
      sigmoid_table_435_2_sva <= sigmoid_table_435_2_sva_dfm_1;
      sigmoid_table_435_5_sva <= sigmoid_table_435_5_sva_dfm_1;
      sigmoid_table_434_5_sva <= sigmoid_table_434_5_sva_dfm_1;
      sigmoid_table_433_1_sva <= sigmoid_table_433_1_sva_dfm_1;
      sigmoid_table_433_5_sva <= sigmoid_table_433_5_sva_dfm_1;
      sigmoid_table_432_5_sva <= sigmoid_table_432_5_sva_dfm_1;
      sigmoid_table_431_5_sva <= sigmoid_table_431_5_sva_dfm_1;
      sigmoid_table_430_1_sva <= sigmoid_table_430_1_sva_dfm_1;
      sigmoid_table_430_6_sva <= sigmoid_table_430_6_sva_dfm_1;
      sigmoid_table_429_0_sva <= sigmoid_table_429_0_sva_dfm_1;
      sigmoid_table_429_3_sva <= sigmoid_table_429_3_sva_dfm_1;
      sigmoid_table_429_6_sva <= sigmoid_table_429_6_sva_dfm_1;
      sigmoid_table_428_3_sva <= sigmoid_table_428_3_sva_dfm_1;
      sigmoid_table_428_6_sva <= sigmoid_table_428_6_sva_dfm_1;
      sigmoid_table_427_1_sva <= sigmoid_table_427_1_sva_dfm_1;
      sigmoid_table_427_6_sva <= sigmoid_table_427_6_sva_dfm_1;
      sigmoid_table_426_0_sva <= sigmoid_table_426_0_sva_dfm_1;
      sigmoid_table_426_6_sva <= sigmoid_table_426_6_sva_dfm_1;
      sigmoid_table_425_6_sva <= sigmoid_table_425_6_sva_dfm_1;
      sigmoid_table_424_1_sva <= sigmoid_table_424_1_sva_dfm_1;
      sigmoid_table_424_6_sva <= sigmoid_table_424_6_sva_dfm_1;
      sigmoid_table_423_2_sva <= sigmoid_table_423_2_sva_dfm_1;
      sigmoid_table_423_6_sva <= sigmoid_table_423_6_sva_dfm_1;
      sigmoid_table_422_6_sva <= sigmoid_table_422_6_sva_dfm_1;
      sigmoid_table_421_0_sva <= sigmoid_table_421_0_sva_dfm_1;
      sigmoid_table_421_6_sva <= sigmoid_table_421_6_sva_dfm_1;
      sigmoid_table_420_6_sva <= sigmoid_table_420_6_sva_dfm_1;
      sigmoid_table_419_6_sva <= sigmoid_table_419_6_sva_dfm_1;
      sigmoid_table_418_0_sva <= sigmoid_table_418_0_sva_dfm_1;
      sigmoid_table_417_2_sva <= sigmoid_table_417_2_sva_dfm_1;
      sigmoid_table_416_3_sva <= sigmoid_table_416_3_sva_dfm_1;
      sigmoid_table_415_3_sva <= sigmoid_table_415_3_sva_dfm_1;
      sigmoid_table_414_1_sva <= sigmoid_table_414_1_sva_dfm_1;
      sigmoid_table_414_4_sva <= sigmoid_table_414_4_sva_dfm_1;
      sigmoid_table_413_0_sva <= sigmoid_table_413_0_sva_dfm_1;
      sigmoid_table_413_4_sva <= sigmoid_table_413_4_sva_dfm_1;
      sigmoid_table_412_4_sva <= sigmoid_table_412_4_sva_dfm_1;
      sigmoid_table_411_0_sva <= sigmoid_table_411_0_sva_dfm_1;
      sigmoid_table_410_2_sva <= sigmoid_table_410_2_sva_dfm_1;
      sigmoid_table_407_1_sva <= sigmoid_table_407_1_sva_dfm_1;
      sigmoid_table_404_0_sva <= sigmoid_table_404_0_sva_dfm_1;
      sigmoid_table_403_2_sva <= sigmoid_table_403_2_sva_dfm_1;
      sigmoid_table_402_0_sva <= sigmoid_table_402_0_sva_dfm_1;
      sigmoid_table_402_3_sva <= sigmoid_table_402_3_sva_dfm_1;
      sigmoid_table_401_3_sva <= sigmoid_table_401_3_sva_dfm_1;
      sigmoid_table_400_0_sva <= sigmoid_table_400_0_sva_dfm_1;
      sigmoid_table_398_0_sva <= sigmoid_table_398_0_sva_dfm_1;
      sigmoid_table_396_0_sva <= sigmoid_table_396_0_sva_dfm_1;
      sigmoid_table_395_2_sva <= sigmoid_table_395_2_sva_dfm_1;
      sigmoid_table_394_0_sva <= sigmoid_table_394_0_sva_dfm_1;
      sigmoid_table_391_1_sva <= sigmoid_table_391_1_sva_dfm_1;
      sigmoid_table_387_0_sva <= sigmoid_table_387_0_sva_dfm_1;
      sigmoid_table_386_2_sva <= sigmoid_table_386_2_sva_dfm_1;
      sigmoid_table_385_0_sva <= sigmoid_table_385_0_sva_dfm_1;
      sigmoid_table_385_3_sva <= sigmoid_table_385_3_sva_dfm_1;
      sigmoid_table_384_3_sva <= sigmoid_table_384_3_sva_dfm_1;
      sigmoid_table_383_3_sva <= sigmoid_table_383_3_sva_dfm_1;
      sigmoid_table_382_1_sva <= sigmoid_table_382_1_sva_dfm_1;
      sigmoid_table_382_4_sva <= sigmoid_table_382_4_sva_dfm_1;
      sigmoid_table_381_4_sva <= sigmoid_table_381_4_sva_dfm_1;
      sigmoid_table_380_0_sva <= sigmoid_table_380_0_sva_dfm_1;
      sigmoid_table_380_4_sva <= sigmoid_table_380_4_sva_dfm_1;
      sigmoid_table_379_4_sva <= sigmoid_table_379_4_sva_dfm_1;
      sigmoid_table_378_4_sva <= sigmoid_table_378_4_sva_dfm_1;
      sigmoid_table_377_1_sva <= sigmoid_table_377_1_sva_dfm_1;
      sigmoid_table_377_5_sva <= sigmoid_table_377_5_sva_dfm_1;
      sigmoid_table_376_2_sva <= sigmoid_table_376_2_sva_dfm_1;
      sigmoid_table_376_5_sva <= sigmoid_table_376_5_sva_dfm_1;
      sigmoid_table_375_0_sva <= sigmoid_table_375_0_sva_dfm_1;
      sigmoid_table_375_5_sva <= sigmoid_table_375_5_sva_dfm_1;
      sigmoid_table_374_5_sva <= sigmoid_table_374_5_sva_dfm_1;
      sigmoid_table_373_5_sva <= sigmoid_table_373_5_sva_dfm_1;
      sigmoid_table_372_0_sva <= sigmoid_table_372_0_sva_dfm_1;
      sigmoid_table_372_5_sva <= sigmoid_table_372_5_sva_dfm_1;
      sigmoid_table_371_5_sva <= sigmoid_table_371_5_sva_dfm_1;
      sigmoid_table_370_5_sva <= sigmoid_table_370_5_sva_dfm_1;
      sigmoid_table_369_0_sva <= sigmoid_table_369_0_sva_dfm_1;
      sigmoid_table_369_5_sva <= sigmoid_table_369_5_sva_dfm_1;
      sigmoid_table_368_5_sva <= sigmoid_table_368_5_sva_dfm_1;
      sigmoid_table_367_5_sva <= sigmoid_table_367_5_sva_dfm_1;
      sigmoid_table_366_1_sva <= sigmoid_table_366_1_sva_dfm_1;
      sigmoid_table_365_2_sva <= sigmoid_table_365_2_sva_dfm_1;
      sigmoid_table_364_2_sva <= sigmoid_table_364_2_sva_dfm_1;
      sigmoid_table_363_3_sva <= sigmoid_table_363_3_sva_dfm_1;
      sigmoid_table_362_3_sva <= sigmoid_table_362_3_sva_dfm_1;
      sigmoid_table_361_3_sva <= sigmoid_table_361_3_sva_dfm_1;
      sigmoid_table_360_0_sva <= sigmoid_table_360_0_sva_dfm_1;
      sigmoid_table_357_0_sva <= sigmoid_table_357_0_sva_dfm_1;
      sigmoid_table_354_0_sva <= sigmoid_table_354_0_sva_dfm_1;
      sigmoid_table_353_1_sva <= sigmoid_table_353_1_sva_dfm_1;
      sigmoid_table_352_2_sva <= sigmoid_table_352_2_sva_dfm_1;
      sigmoid_table_351_2_sva <= sigmoid_table_351_2_sva_dfm_1;
      sigmoid_table_350_0_sva <= sigmoid_table_350_0_sva_dfm_1;
      sigmoid_table_346_0_sva <= sigmoid_table_346_0_sva_dfm_1;
      sigmoid_table_345_1_sva <= sigmoid_table_345_1_sva_dfm_1;
      sigmoid_table_342_0_sva <= sigmoid_table_342_0_sva_dfm_1;
      sigmoid_table_338_0_sva <= sigmoid_table_338_0_sva_dfm_1;
      sigmoid_table_337_1_sva <= sigmoid_table_337_1_sva_dfm_1;
      sigmoid_table_336_2_sva <= sigmoid_table_336_2_sva_dfm_1;
      sigmoid_table_335_2_sva <= sigmoid_table_335_2_sva_dfm_1;
      sigmoid_table_334_0_sva <= sigmoid_table_334_0_sva_dfm_1;
      sigmoid_table_334_3_sva <= sigmoid_table_334_3_sva_dfm_1;
      sigmoid_table_333_3_sva <= sigmoid_table_333_3_sva_dfm_1;
      sigmoid_table_332_3_sva <= sigmoid_table_332_3_sva_dfm_1;
      sigmoid_table_331_3_sva <= sigmoid_table_331_3_sva_dfm_1;
      sigmoid_table_330_3_sva <= sigmoid_table_330_3_sva_dfm_1;
      sigmoid_table_329_0_sva <= sigmoid_table_329_0_sva_dfm_1;
      sigmoid_table_329_4_sva <= sigmoid_table_329_4_sva_dfm_1;
      sigmoid_table_328_1_sva <= sigmoid_table_328_1_sva_dfm_1;
      sigmoid_table_328_4_sva <= sigmoid_table_328_4_sva_dfm_1;
      sigmoid_table_327_4_sva <= sigmoid_table_327_4_sva_dfm_1;
      sigmoid_table_326_4_sva <= sigmoid_table_326_4_sva_dfm_1;
      sigmoid_table_325_4_sva <= sigmoid_table_325_4_sva_dfm_1;
      sigmoid_table_324_0_sva <= sigmoid_table_324_0_sva_dfm_1;
      sigmoid_table_324_4_sva <= sigmoid_table_324_4_sva_dfm_1;
      sigmoid_table_323_4_sva <= sigmoid_table_323_4_sva_dfm_1;
      sigmoid_table_322_4_sva <= sigmoid_table_322_4_sva_dfm_1;
      sigmoid_table_321_4_sva <= sigmoid_table_321_4_sva_dfm_1;
      sigmoid_table_320_4_sva <= sigmoid_table_320_4_sva_dfm_1;
      sigmoid_table_319_0_sva <= sigmoid_table_319_0_sva_dfm_1;
      sigmoid_table_318_0_sva <= sigmoid_table_318_0_sva_dfm_1;
      sigmoid_table_317_1_sva <= sigmoid_table_317_1_sva_dfm_1;
      sigmoid_table_316_2_sva <= sigmoid_table_316_2_sva_dfm_1;
      sigmoid_table_315_2_sva <= sigmoid_table_315_2_sva_dfm_1;
      sigmoid_table_314_2_sva <= sigmoid_table_314_2_sva_dfm_1;
      sigmoid_table_313_0_sva <= sigmoid_table_313_0_sva_dfm_1;
      sigmoid_table_312_0_sva <= sigmoid_table_312_0_sva_dfm_1;
      sigmoid_table_307_0_sva <= sigmoid_table_307_0_sva_dfm_1;
      sigmoid_table_306_0_sva <= sigmoid_table_306_0_sva_dfm_1;
      sigmoid_table_305_1_sva <= sigmoid_table_305_1_sva_dfm_1;
      sigmoid_table_304_1_sva <= sigmoid_table_304_1_sva_dfm_1;
      sigmoid_table_300_0_sva <= sigmoid_table_300_0_sva_dfm_1;
      sigmoid_table_299_0_sva <= sigmoid_table_299_0_sva_dfm_1;
      sigmoid_table_292_0_sva <= sigmoid_table_292_0_sva_dfm_1;
      sigmoid_table_291_0_sva <= sigmoid_table_291_0_sva_dfm_1;
      sigmoid_table_290_1_sva <= sigmoid_table_290_1_sva_dfm_1;
      sigmoid_table_289_1_sva <= sigmoid_table_289_1_sva_dfm_1;
      sigmoid_table_288_1_sva <= sigmoid_table_288_1_sva_dfm_1;
      sigmoid_table_287_2_sva <= sigmoid_table_287_2_sva_dfm_1;
      sigmoid_table_286_2_sva <= sigmoid_table_286_2_sva_dfm_1;
      sigmoid_table_285_2_sva <= sigmoid_table_285_2_sva_dfm_1;
      sigmoid_table_284_2_sva <= sigmoid_table_284_2_sva_dfm_1;
      sigmoid_table_283_0_sva <= sigmoid_table_283_0_sva_dfm_1;
      sigmoid_table_283_3_sva <= sigmoid_table_283_3_sva_dfm_1;
      sigmoid_table_282_0_sva <= sigmoid_table_282_0_sva_dfm_1;
      sigmoid_table_282_3_sva <= sigmoid_table_282_3_sva_dfm_1;
      sigmoid_table_281_3_sva <= sigmoid_table_281_3_sva_dfm_1;
      sigmoid_table_280_3_sva <= sigmoid_table_280_3_sva_dfm_1;
      sigmoid_table_279_3_sva <= sigmoid_table_279_3_sva_dfm_1;
      sigmoid_table_278_3_sva <= sigmoid_table_278_3_sva_dfm_1;
      sigmoid_table_277_3_sva <= sigmoid_table_277_3_sva_dfm_1;
      sigmoid_table_276_3_sva <= sigmoid_table_276_3_sva_dfm_1;
      sigmoid_table_275_3_sva <= sigmoid_table_275_3_sva_dfm_1;
      sigmoid_table_274_3_sva <= sigmoid_table_274_3_sva_dfm_1;
      sigmoid_table_273_0_sva <= sigmoid_table_273_0_sva_dfm_1;
      sigmoid_table_272_0_sva <= sigmoid_table_272_0_sva_dfm_1;
      sigmoid_table_271_0_sva <= sigmoid_table_271_0_sva_dfm_1;
      sigmoid_table_270_1_sva <= sigmoid_table_270_1_sva_dfm_1;
      sigmoid_table_269_1_sva <= sigmoid_table_269_1_sva_dfm_1;
      sigmoid_table_268_1_sva <= sigmoid_table_268_1_sva_dfm_1;
      sigmoid_table_261_0_sva <= sigmoid_table_261_0_sva_dfm_1;
      sigmoid_table_260_0_sva <= sigmoid_table_260_0_sva_dfm_1;
      sigmoid_table_259_0_sva <= sigmoid_table_259_0_sva_dfm_1;
      sigmoid_table_246_0_sva <= sigmoid_table_246_0_sva_dfm_1;
      sigmoid_table_245_0_sva <= sigmoid_table_245_0_sva_dfm_1;
      sigmoid_table_244_0_sva <= sigmoid_table_244_0_sva_dfm_1;
      sigmoid_table_243_0_sva <= sigmoid_table_243_0_sva_dfm_1;
      sigmoid_table_242_1_sva <= sigmoid_table_242_1_sva_dfm_1;
      sigmoid_table_241_1_sva <= sigmoid_table_241_1_sva_dfm_1;
      sigmoid_table_240_1_sva <= sigmoid_table_240_1_sva_dfm_1;
      sigmoid_table_239_1_sva <= sigmoid_table_239_1_sva_dfm_1;
      sigmoid_table_238_2_sva <= sigmoid_table_238_2_sva_dfm_1;
      sigmoid_table_237_2_sva <= sigmoid_table_237_2_sva_dfm_1;
      sigmoid_table_236_2_sva <= sigmoid_table_236_2_sva_dfm_1;
      sigmoid_table_235_2_sva <= sigmoid_table_235_2_sva_dfm_1;
      sigmoid_table_234_2_sva <= sigmoid_table_234_2_sva_dfm_1;
      sigmoid_table_233_2_sva <= sigmoid_table_233_2_sva_dfm_1;
      sigmoid_table_232_2_sva <= sigmoid_table_232_2_sva_dfm_1;
      sigmoid_table_231_2_sva <= sigmoid_table_231_2_sva_dfm_1;
      sigmoid_table_230_2_sva <= sigmoid_table_230_2_sva_dfm_1;
      sigmoid_table_229_2_sva <= sigmoid_table_229_2_sva_dfm_1;
      sigmoid_table_228_0_sva <= sigmoid_table_228_0_sva_dfm_1;
      sigmoid_table_227_0_sva <= sigmoid_table_227_0_sva_dfm_1;
      sigmoid_table_226_0_sva <= sigmoid_table_226_0_sva_dfm_1;
      sigmoid_table_225_0_sva <= sigmoid_table_225_0_sva_dfm_1;
      sigmoid_table_224_0_sva <= sigmoid_table_224_0_sva_dfm_1;
      sigmoid_table_223_0_sva <= sigmoid_table_223_0_sva_dfm_1;
      sigmoid_table_201_0_sva <= sigmoid_table_201_0_sva_dfm_1;
      sigmoid_table_200_0_sva <= sigmoid_table_200_0_sva_dfm_1;
      sigmoid_table_199_0_sva <= sigmoid_table_199_0_sva_dfm_1;
      sigmoid_table_198_0_sva <= sigmoid_table_198_0_sva_dfm_1;
      sigmoid_table_197_0_sva <= sigmoid_table_197_0_sva_dfm_1;
      sigmoid_table_196_0_sva <= sigmoid_table_196_0_sva_dfm_1;
      sigmoid_table_195_0_sva <= sigmoid_table_195_0_sva_dfm_1;
      sigmoid_table_194_0_sva <= sigmoid_table_194_0_sva_dfm_1;
      sigmoid_table_193_1_sva <= sigmoid_table_193_1_sva_dfm_1;
      sigmoid_table_192_1_sva <= sigmoid_table_192_1_sva_dfm_1;
      sigmoid_table_191_1_sva <= sigmoid_table_191_1_sva_dfm_1;
      sigmoid_table_190_1_sva <= sigmoid_table_190_1_sva_dfm_1;
      sigmoid_table_189_1_sva <= sigmoid_table_189_1_sva_dfm_1;
      sigmoid_table_188_1_sva <= sigmoid_table_188_1_sva_dfm_1;
      sigmoid_table_187_1_sva <= sigmoid_table_187_1_sva_dfm_1;
      sigmoid_table_186_1_sva <= sigmoid_table_186_1_sva_dfm_1;
      sigmoid_table_185_1_sva <= sigmoid_table_185_1_sva_dfm_1;
      sigmoid_table_184_1_sva <= sigmoid_table_184_1_sva_dfm_1;
      sigmoid_table_157_0_sva <= sigmoid_table_157_0_sva_dfm_1;
      sigmoid_table_156_0_sva <= sigmoid_table_156_0_sva_dfm_1;
      sigmoid_table_155_0_sva <= sigmoid_table_155_0_sva_dfm_1;
      sigmoid_table_154_0_sva <= sigmoid_table_154_0_sva_dfm_1;
      sigmoid_table_153_0_sva <= sigmoid_table_153_0_sva_dfm_1;
      sigmoid_table_152_0_sva <= sigmoid_table_152_0_sva_dfm_1;
      sigmoid_table_151_0_sva <= sigmoid_table_151_0_sva_dfm_1;
      sigmoid_table_150_0_sva <= sigmoid_table_150_0_sva_dfm_1;
      sigmoid_table_149_0_sva <= sigmoid_table_149_0_sva_dfm_1;
      sigmoid_table_148_0_sva <= sigmoid_table_148_0_sva_dfm_1;
      sigmoid_table_147_0_sva <= sigmoid_table_147_0_sva_dfm_1;
      sigmoid_table_146_0_sva <= sigmoid_table_146_0_sva_dfm_1;
      sigmoid_table_145_0_sva <= sigmoid_table_145_0_sva_dfm_1;
      sigmoid_table_144_0_sva <= sigmoid_table_144_0_sva_dfm_1;
      sigmoid_table_143_0_sva <= sigmoid_table_143_0_sva_dfm_1;
      sigmoid_table_142_0_sva <= sigmoid_table_142_0_sva_dfm_1;
      sigmoid_table_141_0_sva <= sigmoid_table_141_0_sva_dfm_1;
      sigmoid_table_140_0_sva <= sigmoid_table_140_0_sva_dfm_1;
      sigmoid_table_139_0_sva <= sigmoid_table_139_0_sva_dfm_1;
      sigmoid_table_910_0_sva <= sigmoid_table_910_0_sva_dfm_1;
      sigmoid_table_909_0_sva <= sigmoid_table_909_0_sva_dfm_1;
      sigmoid_table_908_0_sva <= sigmoid_table_908_0_sva_dfm_1;
      sigmoid_table_907_0_sva <= sigmoid_table_907_0_sva_dfm_1;
      sigmoid_table_906_0_sva <= sigmoid_table_906_0_sva_dfm_1;
      sigmoid_table_905_0_sva <= sigmoid_table_905_0_sva_dfm_1;
      sigmoid_table_904_0_sva <= sigmoid_table_904_0_sva_dfm_1;
      sigmoid_table_903_0_sva <= sigmoid_table_903_0_sva_dfm_1;
      sigmoid_table_902_0_sva <= sigmoid_table_902_0_sva_dfm_1;
      sigmoid_table_901_0_sva <= sigmoid_table_901_0_sva_dfm_1;
      sigmoid_table_900_0_sva <= sigmoid_table_900_0_sva_dfm_1;
      sigmoid_table_899_0_sva <= sigmoid_table_899_0_sva_dfm_1;
      sigmoid_table_898_0_sva <= sigmoid_table_898_0_sva_dfm_1;
      sigmoid_table_897_0_sva <= sigmoid_table_897_0_sva_dfm_1;
      sigmoid_table_896_0_sva <= sigmoid_table_896_0_sva_dfm_1;
      sigmoid_table_895_0_sva <= sigmoid_table_895_0_sva_dfm_1;
      sigmoid_table_894_0_sva <= sigmoid_table_894_0_sva_dfm_1;
      sigmoid_table_893_0_sva <= sigmoid_table_893_0_sva_dfm_1;
      sigmoid_table_892_0_sva <= sigmoid_table_892_0_sva_dfm_1;
      sigmoid_table_891_0_sva <= sigmoid_table_891_0_sva_dfm_1;
      sigmoid_table_890_0_sva <= sigmoid_table_890_0_sva_dfm_1;
      sigmoid_table_889_0_sva <= sigmoid_table_889_0_sva_dfm_1;
      sigmoid_table_888_0_sva <= sigmoid_table_888_0_sva_dfm_1;
      sigmoid_table_887_0_sva <= sigmoid_table_887_0_sva_dfm_1;
      sigmoid_table_886_0_sva <= sigmoid_table_886_0_sva_dfm_1;
      sigmoid_table_885_0_sva <= sigmoid_table_885_0_sva_dfm_1;
      sigmoid_table_852_1_sva <= sigmoid_table_852_1_sva_dfm_1;
      sigmoid_table_851_1_sva <= sigmoid_table_851_1_sva_dfm_1;
      sigmoid_table_850_1_sva <= sigmoid_table_850_1_sva_dfm_1;
      sigmoid_table_849_1_sva <= sigmoid_table_849_1_sva_dfm_1;
      sigmoid_table_848_1_sva <= sigmoid_table_848_1_sva_dfm_1;
      sigmoid_table_847_1_sva <= sigmoid_table_847_1_sva_dfm_1;
      sigmoid_table_846_1_sva <= sigmoid_table_846_1_sva_dfm_1;
      sigmoid_table_845_1_sva <= sigmoid_table_845_1_sva_dfm_1;
      sigmoid_table_844_1_sva <= sigmoid_table_844_1_sva_dfm_1;
      sigmoid_table_843_1_sva <= sigmoid_table_843_1_sva_dfm_1;
      sigmoid_table_842_1_sva <= sigmoid_table_842_1_sva_dfm_1;
      sigmoid_table_841_1_sva <= sigmoid_table_841_1_sva_dfm_1;
      sigmoid_table_840_0_sva <= sigmoid_table_840_0_sva_dfm_1;
      sigmoid_table_839_0_sva <= sigmoid_table_839_0_sva_dfm_1;
      sigmoid_table_838_0_sva <= sigmoid_table_838_0_sva_dfm_1;
      sigmoid_table_837_0_sva <= sigmoid_table_837_0_sva_dfm_1;
      sigmoid_table_836_0_sva <= sigmoid_table_836_0_sva_dfm_1;
      sigmoid_table_835_0_sva <= sigmoid_table_835_0_sva_dfm_1;
      sigmoid_table_834_0_sva <= sigmoid_table_834_0_sva_dfm_1;
      sigmoid_table_833_0_sva <= sigmoid_table_833_0_sva_dfm_1;
      sigmoid_table_832_0_sva <= sigmoid_table_832_0_sva_dfm_1;
      sigmoid_table_831_0_sva <= sigmoid_table_831_0_sva_dfm_1;
      sigmoid_table_807_0_sva <= sigmoid_table_807_0_sva_dfm_1;
      sigmoid_table_807_2_sva <= sigmoid_table_807_2_sva_dfm_1;
      sigmoid_table_806_0_sva <= sigmoid_table_806_0_sva_dfm_1;
      sigmoid_table_806_2_sva <= sigmoid_table_806_2_sva_dfm_1;
      sigmoid_table_805_0_sva <= sigmoid_table_805_0_sva_dfm_1;
      sigmoid_table_805_2_sva <= sigmoid_table_805_2_sva_dfm_1;
      sigmoid_table_804_0_sva <= sigmoid_table_804_0_sva_dfm_1;
      sigmoid_table_804_2_sva <= sigmoid_table_804_2_sva_dfm_1;
      sigmoid_table_803_0_sva <= sigmoid_table_803_0_sva_dfm_1;
      sigmoid_table_803_2_sva <= sigmoid_table_803_2_sva_dfm_1;
      sigmoid_table_802_0_sva <= sigmoid_table_802_0_sva_dfm_1;
      sigmoid_table_802_2_sva <= sigmoid_table_802_2_sva_dfm_1;
      sigmoid_table_801_2_sva <= sigmoid_table_801_2_sva_dfm_1;
      sigmoid_table_800_2_sva <= sigmoid_table_800_2_sva_dfm_1;
      sigmoid_table_799_2_sva <= sigmoid_table_799_2_sva_dfm_1;
      sigmoid_table_798_2_sva <= sigmoid_table_798_2_sva_dfm_1;
      sigmoid_table_797_2_sva <= sigmoid_table_797_2_sva_dfm_1;
      sigmoid_table_796_2_sva <= sigmoid_table_796_2_sva_dfm_1;
      sigmoid_table_790_1_sva <= sigmoid_table_790_1_sva_dfm_1;
      sigmoid_table_789_1_sva <= sigmoid_table_789_1_sva_dfm_1;
      sigmoid_table_788_1_sva <= sigmoid_table_788_1_sva_dfm_1;
      sigmoid_table_787_1_sva <= sigmoid_table_787_1_sva_dfm_1;
      sigmoid_table_786_1_sva <= sigmoid_table_786_1_sva_dfm_1;
      sigmoid_table_785_0_sva <= sigmoid_table_785_0_sva_dfm_1;
      sigmoid_table_784_0_sva <= sigmoid_table_784_0_sva_dfm_1;
      sigmoid_table_783_0_sva <= sigmoid_table_783_0_sva_dfm_1;
      sigmoid_table_782_0_sva <= sigmoid_table_782_0_sva_dfm_1;
      sigmoid_table_769_0_sva <= sigmoid_table_769_0_sva_dfm_1;
      sigmoid_table_768_0_sva <= sigmoid_table_768_0_sva_dfm_1;
      sigmoid_table_767_0_sva <= sigmoid_table_767_0_sva_dfm_1;
      sigmoid_table_766_0_sva <= sigmoid_table_766_0_sva_dfm_1;
      sigmoid_table_762_3_sva <= sigmoid_table_762_3_sva_dfm_1;
      sigmoid_table_761_3_sva <= sigmoid_table_761_3_sva_dfm_1;
      sigmoid_table_760_3_sva <= sigmoid_table_760_3_sva_dfm_1;
      sigmoid_table_759_1_sva <= sigmoid_table_759_1_sva_dfm_1;
      sigmoid_table_759_3_sva <= sigmoid_table_759_3_sva_dfm_1;
      sigmoid_table_758_1_sva <= sigmoid_table_758_1_sva_dfm_1;
      sigmoid_table_758_3_sva <= sigmoid_table_758_3_sva_dfm_1;
      sigmoid_table_757_1_sva <= sigmoid_table_757_1_sva_dfm_1;
      sigmoid_table_757_3_sva <= sigmoid_table_757_3_sva_dfm_1;
      sigmoid_table_756_0_sva <= sigmoid_table_756_0_sva_dfm_1;
      sigmoid_table_756_3_sva <= sigmoid_table_756_3_sva_dfm_1;
      sigmoid_table_755_0_sva <= sigmoid_table_755_0_sva_dfm_1;
      sigmoid_table_755_3_sva <= sigmoid_table_755_3_sva_dfm_1;
      sigmoid_table_754_0_sva <= sigmoid_table_754_0_sva_dfm_1;
      sigmoid_table_754_3_sva <= sigmoid_table_754_3_sva_dfm_1;
      sigmoid_table_753_3_sva <= sigmoid_table_753_3_sva_dfm_1;
      sigmoid_table_752_3_sva <= sigmoid_table_752_3_sva_dfm_1;
      sigmoid_table_751_3_sva <= sigmoid_table_751_3_sva_dfm_1;
      sigmoid_table_745_0_sva <= sigmoid_table_745_0_sva_dfm_1;
      sigmoid_table_745_2_sva <= sigmoid_table_745_2_sva_dfm_1;
      sigmoid_table_744_0_sva <= sigmoid_table_744_0_sva_dfm_1;
      sigmoid_table_744_2_sva <= sigmoid_table_744_2_sva_dfm_1;
      sigmoid_table_743_0_sva <= sigmoid_table_743_0_sva_dfm_1;
      sigmoid_table_743_2_sva <= sigmoid_table_743_2_sva_dfm_1;
      sigmoid_table_742_2_sva <= sigmoid_table_742_2_sva_dfm_1;
      sigmoid_table_741_2_sva <= sigmoid_table_741_2_sva_dfm_1;
      sigmoid_table_738_1_sva <= sigmoid_table_738_1_sva_dfm_1;
      sigmoid_table_737_1_sva <= sigmoid_table_737_1_sva_dfm_1;
      sigmoid_table_736_0_sva <= sigmoid_table_736_0_sva_dfm_1;
      sigmoid_table_735_0_sva <= sigmoid_table_735_0_sva_dfm_1;
      sigmoid_table_734_0_sva <= sigmoid_table_734_0_sva_dfm_1;
      sigmoid_table_727_0_sva <= sigmoid_table_727_0_sva_dfm_1;
      sigmoid_table_726_0_sva <= sigmoid_table_726_0_sva_dfm_1;
      sigmoid_table_722_1_sva <= sigmoid_table_722_1_sva_dfm_1;
      sigmoid_table_721_1_sva <= sigmoid_table_721_1_sva_dfm_1;
      sigmoid_table_720_0_sva <= sigmoid_table_720_0_sva_dfm_1;
      sigmoid_table_719_0_sva <= sigmoid_table_719_0_sva_dfm_1;
      sigmoid_table_716_4_sva <= sigmoid_table_716_4_sva_dfm_1;
      sigmoid_table_715_4_sva <= sigmoid_table_715_4_sva_dfm_1;
      sigmoid_table_714_4_sva <= sigmoid_table_714_4_sva_dfm_1;
      sigmoid_table_713_0_sva <= sigmoid_table_713_0_sva_dfm_1;
      sigmoid_table_713_2_sva <= sigmoid_table_713_2_sva_dfm_1;
      sigmoid_table_713_4_sva <= sigmoid_table_713_4_sva_dfm_1;
      sigmoid_table_712_2_sva <= sigmoid_table_712_2_sva_dfm_1;
      sigmoid_table_712_4_sva <= sigmoid_table_712_4_sva_dfm_1;
      sigmoid_table_711_2_sva <= sigmoid_table_711_2_sva_dfm_1;
      sigmoid_table_711_4_sva <= sigmoid_table_711_4_sva_dfm_1;
      sigmoid_table_710_4_sva <= sigmoid_table_710_4_sva_dfm_1;
      sigmoid_table_709_1_sva <= sigmoid_table_709_1_sva_dfm_1;
      sigmoid_table_709_4_sva <= sigmoid_table_709_4_sva_dfm_1;
      sigmoid_table_708_1_sva <= sigmoid_table_708_1_sva_dfm_1;
      sigmoid_table_708_4_sva <= sigmoid_table_708_4_sva_dfm_1;
      sigmoid_table_707_0_sva <= sigmoid_table_707_0_sva_dfm_1;
      sigmoid_table_707_4_sva <= sigmoid_table_707_4_sva_dfm_1;
      sigmoid_table_706_4_sva <= sigmoid_table_706_4_sva_dfm_1;
      sigmoid_table_705_4_sva <= sigmoid_table_705_4_sva_dfm_1;
      sigmoid_table_702_0_sva <= sigmoid_table_702_0_sva_dfm_1;
      sigmoid_table_701_0_sva <= sigmoid_table_701_0_sva_dfm_1;
      sigmoid_table_699_3_sva <= sigmoid_table_699_3_sva_dfm_1;
      sigmoid_table_698_1_sva <= sigmoid_table_698_1_sva_dfm_1;
      sigmoid_table_698_3_sva <= sigmoid_table_698_3_sva_dfm_1;
      sigmoid_table_697_1_sva <= sigmoid_table_697_1_sva_dfm_1;
      sigmoid_table_697_3_sva <= sigmoid_table_697_3_sva_dfm_1;
      sigmoid_table_696_0_sva <= sigmoid_table_696_0_sva_dfm_1;
      sigmoid_table_696_3_sva <= sigmoid_table_696_3_sva_dfm_1;
      sigmoid_table_695_3_sva <= sigmoid_table_695_3_sva_dfm_1;
      sigmoid_table_692_0_sva <= sigmoid_table_692_0_sva_dfm_1;
      sigmoid_table_692_2_sva <= sigmoid_table_692_2_sva_dfm_1;
      sigmoid_table_691_0_sva <= sigmoid_table_691_0_sva_dfm_1;
      sigmoid_table_691_2_sva <= sigmoid_table_691_2_sva_dfm_1;
      sigmoid_table_690_2_sva <= sigmoid_table_690_2_sva_dfm_1;
      sigmoid_table_688_1_sva <= sigmoid_table_688_1_sva_dfm_1;
      sigmoid_table_687_0_sva <= sigmoid_table_687_0_sva_dfm_1;
      sigmoid_table_683_0_sva <= sigmoid_table_683_0_sva_dfm_1;
      sigmoid_table_680_1_sva <= sigmoid_table_680_1_sva_dfm_1;
      sigmoid_table_679_0_sva <= sigmoid_table_679_0_sva_dfm_1;
      sigmoid_table_675_0_sva <= sigmoid_table_675_0_sva_dfm_1;
      sigmoid_table_675_2_sva <= sigmoid_table_675_2_sva_dfm_1;
      sigmoid_table_674_2_sva <= sigmoid_table_674_2_sva_dfm_1;
      sigmoid_table_672_1_sva <= sigmoid_table_672_1_sva_dfm_1;
      sigmoid_table_671_0_sva <= sigmoid_table_671_0_sva_dfm_1;
      sigmoid_table_669_5_sva <= sigmoid_table_669_5_sva_dfm_1;
      sigmoid_table_668_0_sva <= sigmoid_table_668_0_sva_dfm_1;
      sigmoid_table_668_5_sva <= sigmoid_table_668_5_sva_dfm_1;
      sigmoid_table_667_5_sva <= sigmoid_table_667_5_sva_dfm_1;
      sigmoid_table_666_3_sva <= sigmoid_table_666_3_sva_dfm_1;
      sigmoid_table_666_5_sva <= sigmoid_table_666_5_sva_dfm_1;
      sigmoid_table_665_1_sva <= sigmoid_table_665_1_sva_dfm_1;
      sigmoid_table_665_3_sva <= sigmoid_table_665_3_sva_dfm_1;
      sigmoid_table_665_5_sva <= sigmoid_table_665_5_sva_dfm_1;
      sigmoid_table_664_3_sva <= sigmoid_table_664_3_sva_dfm_1;
      sigmoid_table_664_5_sva <= sigmoid_table_664_5_sva_dfm_1;
      sigmoid_table_663_5_sva <= sigmoid_table_663_5_sva_dfm_1;
      sigmoid_table_662_5_sva <= sigmoid_table_662_5_sva_dfm_1;
      sigmoid_table_661_0_sva <= sigmoid_table_661_0_sva_dfm_1;
      sigmoid_table_661_2_sva <= sigmoid_table_661_2_sva_dfm_1;
      sigmoid_table_661_5_sva <= sigmoid_table_661_5_sva_dfm_1;
      sigmoid_table_660_5_sva <= sigmoid_table_660_5_sva_dfm_1;
      sigmoid_table_659_1_sva <= sigmoid_table_659_1_sva_dfm_1;
      sigmoid_table_659_5_sva <= sigmoid_table_659_5_sva_dfm_1;
      sigmoid_table_658_0_sva <= sigmoid_table_658_0_sva_dfm_1;
      sigmoid_table_658_5_sva <= sigmoid_table_658_5_sva_dfm_1;
      sigmoid_table_653_1_sva <= sigmoid_table_653_1_sva_dfm_1;
      sigmoid_table_651_4_sva <= sigmoid_table_651_4_sva_dfm_1;
      sigmoid_table_650_0_sva <= sigmoid_table_650_0_sva_dfm_1;
      sigmoid_table_650_2_sva <= sigmoid_table_650_2_sva_dfm_1;
      sigmoid_table_650_4_sva <= sigmoid_table_650_4_sva_dfm_1;
      sigmoid_table_649_2_sva <= sigmoid_table_649_2_sva_dfm_1;
      sigmoid_table_649_4_sva <= sigmoid_table_649_4_sva_dfm_1;
      sigmoid_table_648_1_sva <= sigmoid_table_648_1_sva_dfm_1;
      sigmoid_table_648_4_sva <= sigmoid_table_648_4_sva_dfm_1;
      sigmoid_table_647_0_sva <= sigmoid_table_647_0_sva_dfm_1;
      sigmoid_table_647_4_sva <= sigmoid_table_647_4_sva_dfm_1;
      sigmoid_table_643_1_sva <= sigmoid_table_643_1_sva_dfm_1;
      sigmoid_table_643_3_sva <= sigmoid_table_643_3_sva_dfm_1;
      sigmoid_table_642_0_sva <= sigmoid_table_642_0_sva_dfm_1;
      sigmoid_table_642_3_sva <= sigmoid_table_642_3_sva_dfm_1;
      sigmoid_table_640_0_sva <= sigmoid_table_640_0_sva_dfm_1;
      sigmoid_table_640_2_sva <= sigmoid_table_640_2_sva_dfm_1;
      sigmoid_table_639_2_sva <= sigmoid_table_639_2_sva_dfm_1;
      sigmoid_table_638_1_sva <= sigmoid_table_638_1_sva_dfm_1;
      sigmoid_table_635_0_sva <= sigmoid_table_635_0_sva_dfm_1;
      sigmoid_table_633_0_sva <= sigmoid_table_633_0_sva_dfm_1;
      sigmoid_table_631_0_sva <= sigmoid_table_631_0_sva_dfm_1;
      sigmoid_table_631_2_sva <= sigmoid_table_631_2_sva_dfm_1;
      sigmoid_table_630_2_sva <= sigmoid_table_630_2_sva_dfm_1;
      sigmoid_table_629_1_sva <= sigmoid_table_629_1_sva_dfm_1;
      sigmoid_table_625_1_sva <= sigmoid_table_625_1_sva_dfm_1;
      sigmoid_table_625_3_sva <= sigmoid_table_625_3_sva_dfm_1;
      sigmoid_table_624_3_sva <= sigmoid_table_624_3_sva_dfm_1;
      sigmoid_table_622_2_sva <= sigmoid_table_622_2_sva_dfm_1;
      sigmoid_table_621_1_sva <= sigmoid_table_621_1_sva_dfm_1;
      sigmoid_table_619_6_sva <= sigmoid_table_619_6_sva_dfm_1;
      sigmoid_table_618_6_sva <= sigmoid_table_618_6_sva_dfm_1;
      sigmoid_table_617_0_sva <= sigmoid_table_617_0_sva_dfm_1;
      sigmoid_table_617_6_sva <= sigmoid_table_617_6_sva_dfm_1;
      sigmoid_table_616_4_sva <= sigmoid_table_616_4_sva_dfm_1;
      sigmoid_table_616_6_sva <= sigmoid_table_616_6_sva_dfm_1;
      sigmoid_table_615_0_sva <= sigmoid_table_615_0_sva_dfm_1;
      sigmoid_table_615_2_sva <= sigmoid_table_615_2_sva_dfm_1;
      sigmoid_table_615_4_sva <= sigmoid_table_615_4_sva_dfm_1;
      sigmoid_table_615_6_sva <= sigmoid_table_615_6_sva_dfm_1;
      sigmoid_table_614_4_sva <= sigmoid_table_614_4_sva_dfm_1;
      sigmoid_table_614_6_sva <= sigmoid_table_614_6_sva_dfm_1;
      sigmoid_table_613_4_sva <= sigmoid_table_613_4_sva_dfm_1;
      sigmoid_table_613_6_sva <= sigmoid_table_613_6_sva_dfm_1;
      sigmoid_table_612_6_sva <= sigmoid_table_612_6_sva_dfm_1;
      sigmoid_table_611_6_sva <= sigmoid_table_611_6_sva_dfm_1;
      sigmoid_table_610_0_sva <= sigmoid_table_610_0_sva_dfm_1;
      sigmoid_table_610_3_sva <= sigmoid_table_610_3_sva_dfm_1;
      sigmoid_table_610_6_sva <= sigmoid_table_610_6_sva_dfm_1;
      sigmoid_table_609_6_sva <= sigmoid_table_609_6_sva_dfm_1;
      sigmoid_table_608_0_sva <= sigmoid_table_608_0_sva_dfm_1;
      sigmoid_table_608_2_sva <= sigmoid_table_608_2_sva_dfm_1;
      sigmoid_table_608_6_sva <= sigmoid_table_608_6_sva_dfm_1;
      sigmoid_table_607_1_sva <= sigmoid_table_607_1_sva_dfm_1;
      sigmoid_table_607_6_sva <= sigmoid_table_607_6_sva_dfm_1;
      sigmoid_table_606_6_sva <= sigmoid_table_606_6_sva_dfm_1;
      sigmoid_table_605_0_sva <= sigmoid_table_605_0_sva_dfm_1;
      sigmoid_table_600_0_sva <= sigmoid_table_600_0_sva_dfm_1;
      sigmoid_table_599_5_sva <= sigmoid_table_599_5_sva_dfm_1;
      sigmoid_table_598_5_sva <= sigmoid_table_598_5_sva_dfm_1;
      sigmoid_table_597_0_sva <= sigmoid_table_597_0_sva_dfm_1;
      sigmoid_table_597_3_sva <= sigmoid_table_597_3_sva_dfm_1;
      sigmoid_table_597_5_sva <= sigmoid_table_597_5_sva_dfm_1;
      sigmoid_table_596_5_sva <= sigmoid_table_596_5_sva_dfm_1;
      sigmoid_table_595_2_sva <= sigmoid_table_595_2_sva_dfm_1;
      sigmoid_table_595_5_sva <= sigmoid_table_595_5_sva_dfm_1;
      sigmoid_table_594_0_sva <= sigmoid_table_594_0_sva_dfm_1;
      sigmoid_table_594_5_sva <= sigmoid_table_594_5_sva_dfm_1;
      sigmoid_table_591_0_sva <= sigmoid_table_591_0_sva_dfm_1;
      sigmoid_table_590_4_sva <= sigmoid_table_590_4_sva_dfm_1;
      sigmoid_table_589_4_sva <= sigmoid_table_589_4_sva_dfm_1;
      sigmoid_table_588_4_sva <= sigmoid_table_588_4_sva_dfm_1;
      sigmoid_table_587_0_sva <= sigmoid_table_587_0_sva_dfm_1;
      sigmoid_table_586_1_sva <= sigmoid_table_586_1_sva_dfm_1;
      sigmoid_table_586_3_sva <= sigmoid_table_586_3_sva_dfm_1;
      sigmoid_table_584_0_sva <= sigmoid_table_584_0_sva_dfm_1;
      sigmoid_table_584_2_sva <= sigmoid_table_584_2_sva_dfm_1;
      sigmoid_table_583_1_sva <= sigmoid_table_583_1_sva_dfm_1;
      sigmoid_table_582_9_sva <= sigmoid_table_582_9_sva_dfm_1;
      sigmoid_table_581_9_sva <= sigmoid_table_581_9_sva_dfm_1;
      sigmoid_table_580_0_sva <= sigmoid_table_580_0_sva_dfm_1;
      sigmoid_table_580_9_sva <= sigmoid_table_580_9_sva_dfm_1;
      sigmoid_table_579_0_sva <= sigmoid_table_579_0_sva_dfm_1;
      sigmoid_table_579_2_sva <= sigmoid_table_579_2_sva_dfm_1;
      sigmoid_table_579_9_sva <= sigmoid_table_579_9_sva_dfm_1;
      sigmoid_table_578_1_sva <= sigmoid_table_578_1_sva_dfm_1;
      sigmoid_table_578_9_sva <= sigmoid_table_578_9_sva_dfm_1;
      sigmoid_table_577_9_sva <= sigmoid_table_577_9_sva_dfm_1;
      sigmoid_table_576_9_sva <= sigmoid_table_576_9_sva_dfm_1;
      sigmoid_table_575_0_sva <= sigmoid_table_575_0_sva_dfm_1;
      sigmoid_table_575_3_sva <= sigmoid_table_575_3_sva_dfm_1;
      sigmoid_table_575_9_sva <= sigmoid_table_575_9_sva_dfm_1;
      sigmoid_table_574_9_sva <= sigmoid_table_574_9_sva_dfm_1;
      sigmoid_table_573_9_sva <= sigmoid_table_573_9_sva_dfm_1;
      sigmoid_table_572_9_sva <= sigmoid_table_572_9_sva_dfm_1;
      sigmoid_table_571_9_sva <= sigmoid_table_571_9_sva_dfm_1;
      sigmoid_table_570_0_sva <= sigmoid_table_570_0_sva_dfm_1;
      sigmoid_table_570_9_sva <= sigmoid_table_570_9_sva_dfm_1;
      sigmoid_table_569_4_sva <= sigmoid_table_569_4_sva_dfm_1;
      sigmoid_table_569_9_sva <= sigmoid_table_569_9_sva_dfm_1;
      sigmoid_table_568_1_sva <= sigmoid_table_568_1_sva_dfm_1;
      sigmoid_table_568_4_sva <= sigmoid_table_568_4_sva_dfm_1;
      sigmoid_table_568_9_sva <= sigmoid_table_568_9_sva_dfm_1;
      sigmoid_table_567_9_sva <= sigmoid_table_567_9_sva_dfm_1;
      sigmoid_table_566_9_sva <= sigmoid_table_566_9_sva_dfm_1;
      sigmoid_table_565_3_sva <= sigmoid_table_565_3_sva_dfm_1;
      sigmoid_table_565_9_sva <= sigmoid_table_565_9_sva_dfm_1;
      sigmoid_table_564_0_sva <= sigmoid_table_564_0_sva_dfm_1;
      sigmoid_table_564_2_sva <= sigmoid_table_564_2_sva_dfm_1;
      sigmoid_table_564_9_sva <= sigmoid_table_564_9_sva_dfm_1;
      sigmoid_table_563_0_sva <= sigmoid_table_563_0_sva_dfm_1;
      sigmoid_table_563_9_sva <= sigmoid_table_563_9_sva_dfm_1;
      sigmoid_table_562_7_sva <= sigmoid_table_562_7_sva_dfm_1;
      sigmoid_table_562_9_sva <= sigmoid_table_562_9_sva_dfm_1;
      sigmoid_table_561_1_sva <= sigmoid_table_561_1_sva_dfm_1;
      sigmoid_table_561_7_sva <= sigmoid_table_561_7_sva_dfm_1;
      sigmoid_table_561_9_sva <= sigmoid_table_561_9_sva_dfm_1;
      sigmoid_table_560_7_sva <= sigmoid_table_560_7_sva_dfm_1;
      sigmoid_table_560_9_sva <= sigmoid_table_560_9_sva_dfm_1;
      sigmoid_table_559_7_sva <= sigmoid_table_559_7_sva_dfm_1;
      sigmoid_table_559_9_sva <= sigmoid_table_559_9_sva_dfm_1;
      sigmoid_table_558_7_sva <= sigmoid_table_558_7_sva_dfm_1;
      sigmoid_table_558_9_sva <= sigmoid_table_558_9_sva_dfm_1;
      sigmoid_table_557_5_sva <= sigmoid_table_557_5_sva_dfm_1;
      sigmoid_table_557_7_sva <= sigmoid_table_557_7_sva_dfm_1;
      sigmoid_table_557_9_sva <= sigmoid_table_557_9_sva_dfm_1;
      sigmoid_table_556_0_sva <= sigmoid_table_556_0_sva_dfm_1;
      sigmoid_table_556_3_sva <= sigmoid_table_556_3_sva_dfm_1;
      sigmoid_table_556_5_sva <= sigmoid_table_556_5_sva_dfm_1;
      sigmoid_table_556_7_sva <= sigmoid_table_556_7_sva_dfm_1;
      sigmoid_table_556_9_sva <= sigmoid_table_556_9_sva_dfm_1;
      sigmoid_table_555_0_sva <= sigmoid_table_555_0_sva_dfm_1;
      sigmoid_table_555_2_sva <= sigmoid_table_555_2_sva_dfm_1;
      sigmoid_table_555_5_sva <= sigmoid_table_555_5_sva_dfm_1;
      sigmoid_table_555_7_sva <= sigmoid_table_555_7_sva_dfm_1;
      sigmoid_table_555_9_sva <= sigmoid_table_555_9_sva_dfm_1;
      sigmoid_table_554_1_sva <= sigmoid_table_554_1_sva_dfm_1;
      sigmoid_table_554_5_sva <= sigmoid_table_554_5_sva_dfm_1;
      sigmoid_table_554_7_sva <= sigmoid_table_554_7_sva_dfm_1;
      sigmoid_table_554_9_sva <= sigmoid_table_554_9_sva_dfm_1;
      sigmoid_table_553_7_sva <= sigmoid_table_553_7_sva_dfm_1;
      sigmoid_table_553_9_sva <= sigmoid_table_553_9_sva_dfm_1;
      sigmoid_table_552_1_sva <= sigmoid_table_552_1_sva_dfm_1;
      sigmoid_table_552_7_sva <= sigmoid_table_552_7_sva_dfm_1;
      sigmoid_table_552_9_sva <= sigmoid_table_552_9_sva_dfm_1;
      sigmoid_table_551_4_sva <= sigmoid_table_551_4_sva_dfm_1;
      sigmoid_table_551_7_sva <= sigmoid_table_551_7_sva_dfm_1;
      sigmoid_table_551_9_sva <= sigmoid_table_551_9_sva_dfm_1;
      sigmoid_table_550_4_sva <= sigmoid_table_550_4_sva_dfm_1;
      sigmoid_table_550_7_sva <= sigmoid_table_550_7_sva_dfm_1;
      sigmoid_table_550_9_sva <= sigmoid_table_550_9_sva_dfm_1;
      sigmoid_table_549_4_sva <= sigmoid_table_549_4_sva_dfm_1;
      sigmoid_table_549_7_sva <= sigmoid_table_549_7_sva_dfm_1;
      sigmoid_table_549_9_sva <= sigmoid_table_549_9_sva_dfm_1;
      sigmoid_table_548_7_sva <= sigmoid_table_548_7_sva_dfm_1;
      sigmoid_table_548_9_sva <= sigmoid_table_548_9_sva_dfm_1;
      sigmoid_table_547_3_sva <= sigmoid_table_547_3_sva_dfm_1;
      sigmoid_table_547_7_sva <= sigmoid_table_547_7_sva_dfm_1;
      sigmoid_table_547_9_sva <= sigmoid_table_547_9_sva_dfm_1;
      sigmoid_table_546_2_sva <= sigmoid_table_546_2_sva_dfm_1;
      sigmoid_table_546_7_sva <= sigmoid_table_546_7_sva_dfm_1;
      sigmoid_table_546_9_sva <= sigmoid_table_546_9_sva_dfm_1;
      sigmoid_table_545_0_sva <= sigmoid_table_545_0_sva_dfm_1;
      sigmoid_table_545_7_sva <= sigmoid_table_545_7_sva_dfm_1;
      sigmoid_table_545_9_sva <= sigmoid_table_545_9_sva_dfm_1;
      sigmoid_table_544_0_sva <= sigmoid_table_544_0_sva_dfm_1;
      sigmoid_table_544_9_sva <= sigmoid_table_544_9_sva_dfm_1;
      sigmoid_table_543_0_sva <= sigmoid_table_543_0_sva_dfm_1;
      sigmoid_table_543_9_sva <= sigmoid_table_543_9_sva_dfm_1;
      sigmoid_table_542_0_sva <= sigmoid_table_542_0_sva_dfm_1;
      sigmoid_table_542_2_sva <= sigmoid_table_542_2_sva_dfm_1;
      sigmoid_table_542_9_sva <= sigmoid_table_542_9_sva_dfm_1;
      sigmoid_table_541_1_sva <= sigmoid_table_541_1_sva_dfm_1;
      sigmoid_table_541_9_sva <= sigmoid_table_541_9_sva_dfm_1;
      sigmoid_table_540_9_sva <= sigmoid_table_540_9_sva_dfm_1;
      sigmoid_table_539_1_sva <= sigmoid_table_539_1_sva_dfm_1;
      sigmoid_table_539_3_sva <= sigmoid_table_539_3_sva_dfm_1;
      sigmoid_table_539_9_sva <= sigmoid_table_539_9_sva_dfm_1;
      sigmoid_table_538_9_sva <= sigmoid_table_538_9_sva_dfm_1;
      sigmoid_table_537_1_sva <= sigmoid_table_537_1_sva_dfm_1;
      sigmoid_table_537_9_sva <= sigmoid_table_537_9_sva_dfm_1;
      sigmoid_table_536_6_sva <= sigmoid_table_536_6_sva_dfm_1;
      sigmoid_table_536_9_sva <= sigmoid_table_536_9_sva_dfm_1;
      sigmoid_table_535_6_sva <= sigmoid_table_535_6_sva_dfm_1;
      sigmoid_table_535_9_sva <= sigmoid_table_535_9_sva_dfm_1;
      sigmoid_table_534_4_sva <= sigmoid_table_534_4_sva_dfm_1;
      sigmoid_table_534_6_sva <= sigmoid_table_534_6_sva_dfm_1;
      sigmoid_table_534_9_sva <= sigmoid_table_534_9_sva_dfm_1;
      sigmoid_table_533_4_sva <= sigmoid_table_533_4_sva_dfm_1;
      sigmoid_table_533_6_sva <= sigmoid_table_533_6_sva_dfm_1;
      sigmoid_table_533_9_sva <= sigmoid_table_533_9_sva_dfm_1;
      sigmoid_table_532_6_sva <= sigmoid_table_532_6_sva_dfm_1;
      sigmoid_table_532_9_sva <= sigmoid_table_532_9_sva_dfm_1;
      sigmoid_table_531_3_sva <= sigmoid_table_531_3_sva_dfm_1;
      sigmoid_table_531_6_sva <= sigmoid_table_531_6_sva_dfm_1;
      sigmoid_table_531_9_sva <= sigmoid_table_531_9_sva_dfm_1;
      sigmoid_table_530_6_sva <= sigmoid_table_530_6_sva_dfm_1;
      sigmoid_table_530_9_sva <= sigmoid_table_530_9_sva_dfm_1;
      sigmoid_table_529_6_sva <= sigmoid_table_529_6_sva_dfm_1;
      sigmoid_table_529_9_sva <= sigmoid_table_529_9_sva_dfm_1;
      sigmoid_table_528_9_sva <= sigmoid_table_528_9_sva_dfm_1;
      sigmoid_table_527_9_sva <= sigmoid_table_527_9_sva_dfm_1;
      sigmoid_table_526_9_sva <= sigmoid_table_526_9_sva_dfm_1;
      sigmoid_table_525_9_sva <= sigmoid_table_525_9_sva_dfm_1;
      sigmoid_table_524_5_sva <= sigmoid_table_524_5_sva_dfm_1;
      sigmoid_table_524_9_sva <= sigmoid_table_524_9_sva_dfm_1;
      sigmoid_table_523_3_sva <= sigmoid_table_523_3_sva_dfm_1;
      sigmoid_table_523_5_sva <= sigmoid_table_523_5_sva_dfm_1;
      sigmoid_table_523_9_sva <= sigmoid_table_523_9_sva_dfm_1;
      sigmoid_table_522_5_sva <= sigmoid_table_522_5_sva_dfm_1;
      sigmoid_table_522_9_sva <= sigmoid_table_522_9_sva_dfm_1;
      sigmoid_table_521_5_sva <= sigmoid_table_521_5_sva_dfm_1;
      sigmoid_table_521_9_sva <= sigmoid_table_521_9_sva_dfm_1;
      sigmoid_table_520_9_sva <= sigmoid_table_520_9_sva_dfm_1;
      sigmoid_table_519_9_sva <= sigmoid_table_519_9_sva_dfm_1;
      sigmoid_table_518_4_sva <= sigmoid_table_518_4_sva_dfm_1;
      sigmoid_table_518_9_sva <= sigmoid_table_518_9_sva_dfm_1;
      sigmoid_table_517_4_sva <= sigmoid_table_517_4_sva_dfm_1;
      sigmoid_table_517_9_sva <= sigmoid_table_517_9_sva_dfm_1;
      sigmoid_table_516_9_sva <= sigmoid_table_516_9_sva_dfm_1;
      sigmoid_table_515_9_sva <= sigmoid_table_515_9_sva_dfm_1;
      sigmoid_table_514_3_sva <= sigmoid_table_514_3_sva_dfm_1;
      sigmoid_table_514_9_sva <= sigmoid_table_514_9_sva_dfm_1;
      sigmoid_table_513_2_sva <= sigmoid_table_513_2_sva_dfm_1;
      sigmoid_table_513_9_sva <= sigmoid_table_513_9_sva_dfm_1;
      sigmoid_table_512_9_sva <= sigmoid_table_512_9_sva_dfm_1;
      sigmoid_table_509_2_sva <= sigmoid_table_509_2_sva_dfm_1;
      sigmoid_table_506_3_sva <= sigmoid_table_506_3_sva_dfm_1;
      sigmoid_table_505_2_sva <= sigmoid_table_505_2_sva_dfm_1;
      sigmoid_table_501_2_sva <= sigmoid_table_501_2_sva_dfm_1;
      sigmoid_table_501_4_sva <= sigmoid_table_501_4_sva_dfm_1;
      sigmoid_table_500_4_sva <= sigmoid_table_500_4_sva_dfm_1;
      sigmoid_table_498_3_sva <= sigmoid_table_498_3_sva_dfm_1;
      sigmoid_table_497_2_sva <= sigmoid_table_497_2_sva_dfm_1;
      sigmoid_table_493_2_sva <= sigmoid_table_493_2_sva_dfm_1;
      sigmoid_table_491_5_sva <= sigmoid_table_491_5_sva_dfm_1;
      sigmoid_table_490_3_sva <= sigmoid_table_490_3_sva_dfm_1;
      sigmoid_table_490_5_sva <= sigmoid_table_490_5_sva_dfm_1;
      sigmoid_table_489_2_sva <= sigmoid_table_489_2_sva_dfm_1;
      sigmoid_table_489_5_sva <= sigmoid_table_489_5_sva_dfm_1;
      sigmoid_table_488_0_sva <= sigmoid_table_488_0_sva_dfm_1;
      sigmoid_table_488_5_sva <= sigmoid_table_488_5_sva_dfm_1;
      sigmoid_table_487_0_sva <= sigmoid_table_487_0_sva_dfm_1;
      sigmoid_table_486_0_sva <= sigmoid_table_486_0_sva_dfm_1;
      sigmoid_table_485_0_sva <= sigmoid_table_485_0_sva_dfm_1;
      sigmoid_table_485_2_sva <= sigmoid_table_485_2_sva_dfm_1;
      sigmoid_table_485_4_sva <= sigmoid_table_485_4_sva_dfm_1;
      sigmoid_table_484_0_sva <= sigmoid_table_484_0_sva_dfm_1;
      sigmoid_table_484_4_sva <= sigmoid_table_484_4_sva_dfm_1;
      sigmoid_table_483_0_sva <= sigmoid_table_483_0_sva_dfm_1;
      sigmoid_table_482_1_sva <= sigmoid_table_482_1_sva_dfm_1;
      sigmoid_table_482_3_sva <= sigmoid_table_482_3_sva_dfm_1;
      sigmoid_table_480_1_sva <= sigmoid_table_480_1_sva_dfm_1;
      sigmoid_table_479_8_sva <= sigmoid_table_479_8_sva_dfm_1;
      sigmoid_table_478_8_sva <= sigmoid_table_478_8_sva_dfm_1;
      sigmoid_table_477_8_sva <= sigmoid_table_477_8_sva_dfm_1;
      sigmoid_table_476_8_sva <= sigmoid_table_476_8_sva_dfm_1;
      sigmoid_table_475_8_sva <= sigmoid_table_475_8_sva_dfm_1;
      sigmoid_table_474_8_sva <= sigmoid_table_474_8_sva_dfm_1;
      sigmoid_table_473_3_sva <= sigmoid_table_473_3_sva_dfm_1;
      sigmoid_table_473_8_sva <= sigmoid_table_473_8_sva_dfm_1;
      sigmoid_table_472_0_sva <= sigmoid_table_472_0_sva_dfm_1;
      sigmoid_table_472_2_sva <= sigmoid_table_472_2_sva_dfm_1;
      sigmoid_table_472_8_sva <= sigmoid_table_472_8_sva_dfm_1;
      sigmoid_table_471_0_sva <= sigmoid_table_471_0_sva_dfm_1;
      sigmoid_table_471_8_sva <= sigmoid_table_471_8_sva_dfm_1;
      sigmoid_table_470_0_sva <= sigmoid_table_470_0_sva_dfm_1;
      sigmoid_table_470_6_sva <= sigmoid_table_470_6_sva_dfm_1;
      sigmoid_table_470_8_sva <= sigmoid_table_470_8_sva_dfm_1;
      sigmoid_table_469_1_sva <= sigmoid_table_469_1_sva_dfm_1;
      sigmoid_table_469_6_sva <= sigmoid_table_469_6_sva_dfm_1;
      sigmoid_table_469_8_sva <= sigmoid_table_469_8_sva_dfm_1;
      sigmoid_table_468_4_sva <= sigmoid_table_468_4_sva_dfm_1;
      sigmoid_table_468_6_sva <= sigmoid_table_468_6_sva_dfm_1;
      sigmoid_table_468_8_sva <= sigmoid_table_468_8_sva_dfm_1;
      sigmoid_table_467_4_sva <= sigmoid_table_467_4_sva_dfm_1;
      sigmoid_table_467_6_sva <= sigmoid_table_467_6_sva_dfm_1;
      sigmoid_table_467_8_sva <= sigmoid_table_467_8_sva_dfm_1;
      sigmoid_table_466_6_sva <= sigmoid_table_466_6_sva_dfm_1;
      sigmoid_table_466_8_sva <= sigmoid_table_466_8_sva_dfm_1;
      sigmoid_table_465_6_sva <= sigmoid_table_465_6_sva_dfm_1;
      sigmoid_table_465_8_sva <= sigmoid_table_465_8_sva_dfm_1;
      sigmoid_table_464_3_sva <= sigmoid_table_464_3_sva_dfm_1;
      sigmoid_table_464_6_sva <= sigmoid_table_464_6_sva_dfm_1;
      sigmoid_table_464_8_sva <= sigmoid_table_464_8_sva_dfm_1;
      sigmoid_table_463_0_sva <= sigmoid_table_463_0_sva_dfm_1;
      sigmoid_table_463_2_sva <= sigmoid_table_463_2_sva_dfm_1;
      sigmoid_table_463_6_sva <= sigmoid_table_463_6_sva_dfm_1;
      sigmoid_table_463_8_sva <= sigmoid_table_463_8_sva_dfm_1;
      sigmoid_table_462_0_sva <= sigmoid_table_462_0_sva_dfm_1;
      sigmoid_table_462_6_sva <= sigmoid_table_462_6_sva_dfm_1;
      sigmoid_table_462_8_sva <= sigmoid_table_462_8_sva_dfm_1;
      sigmoid_table_461_8_sva <= sigmoid_table_461_8_sva_dfm_1;
      sigmoid_table_460_1_sva <= sigmoid_table_460_1_sva_dfm_1;
      sigmoid_table_460_8_sva <= sigmoid_table_460_8_sva_dfm_1;
      sigmoid_table_459_8_sva <= sigmoid_table_459_8_sva_dfm_1;
      sigmoid_table_458_8_sva <= sigmoid_table_458_8_sva_dfm_1;
      sigmoid_table_457_8_sva <= sigmoid_table_457_8_sva_dfm_1;
      sigmoid_table_456_0_sva <= sigmoid_table_456_0_sva_dfm_1;
      sigmoid_table_456_5_sva <= sigmoid_table_456_5_sva_dfm_1;
      sigmoid_table_456_8_sva <= sigmoid_table_456_8_sva_dfm_1;
      sigmoid_table_455_0_sva <= sigmoid_table_455_0_sva_dfm_1;
      sigmoid_table_455_3_sva <= sigmoid_table_455_3_sva_dfm_1;
      sigmoid_table_455_5_sva <= sigmoid_table_455_5_sva_dfm_1;
      sigmoid_table_455_8_sva <= sigmoid_table_455_8_sva_dfm_1;
      sigmoid_table_454_5_sva <= sigmoid_table_454_5_sva_dfm_1;
      sigmoid_table_454_8_sva <= sigmoid_table_454_8_sva_dfm_1;
      sigmoid_table_453_5_sva <= sigmoid_table_453_5_sva_dfm_1;
      sigmoid_table_453_8_sva <= sigmoid_table_453_8_sva_dfm_1;
      sigmoid_table_452_5_sva <= sigmoid_table_452_5_sva_dfm_1;
      sigmoid_table_452_8_sva <= sigmoid_table_452_8_sva_dfm_1;
      sigmoid_table_451_8_sva <= sigmoid_table_451_8_sva_dfm_1;
      sigmoid_table_450_0_sva <= sigmoid_table_450_0_sva_dfm_1;
      sigmoid_table_450_8_sva <= sigmoid_table_450_8_sva_dfm_1;
      sigmoid_table_449_4_sva <= sigmoid_table_449_4_sva_dfm_1;
      sigmoid_table_449_8_sva <= sigmoid_table_449_8_sva_dfm_1;
      sigmoid_table_448_4_sva <= sigmoid_table_448_4_sva_dfm_1;
      sigmoid_table_448_8_sva <= sigmoid_table_448_8_sva_dfm_1;
      sigmoid_table_447_4_sva <= sigmoid_table_447_4_sva_dfm_1;
      sigmoid_table_447_8_sva <= sigmoid_table_447_8_sva_dfm_1;
      sigmoid_table_446_0_sva <= sigmoid_table_446_0_sva_dfm_1;
      sigmoid_table_446_8_sva <= sigmoid_table_446_8_sva_dfm_1;
      sigmoid_table_445_1_sva <= sigmoid_table_445_1_sva_dfm_1;
      sigmoid_table_445_3_sva <= sigmoid_table_445_3_sva_dfm_1;
      sigmoid_table_445_8_sva <= sigmoid_table_445_8_sva_dfm_1;
      sigmoid_table_444_8_sva <= sigmoid_table_444_8_sva_dfm_1;
      sigmoid_table_443_8_sva <= sigmoid_table_443_8_sva_dfm_1;
      sigmoid_table_442_8_sva <= sigmoid_table_442_8_sva_dfm_1;
      sigmoid_table_441_0_sva <= sigmoid_table_441_0_sva_dfm_1;
      sigmoid_table_440_1_sva <= sigmoid_table_440_1_sva_dfm_1;
      sigmoid_table_438_0_sva <= sigmoid_table_438_0_sva_dfm_1;
      sigmoid_table_438_2_sva <= sigmoid_table_438_2_sva_dfm_1;
      sigmoid_table_437_1_sva <= sigmoid_table_437_1_sva_dfm_1;
      sigmoid_table_434_0_sva <= sigmoid_table_434_0_sva_dfm_1;
      sigmoid_table_434_3_sva <= sigmoid_table_434_3_sva_dfm_1;
      sigmoid_table_432_2_sva <= sigmoid_table_432_2_sva_dfm_1;
      sigmoid_table_431_0_sva <= sigmoid_table_431_0_sva_dfm_1;
      sigmoid_table_428_0_sva <= sigmoid_table_428_0_sva_dfm_1;
      sigmoid_table_427_4_sva <= sigmoid_table_427_4_sva_dfm_1;
      sigmoid_table_426_4_sva <= sigmoid_table_426_4_sva_dfm_1;
      sigmoid_table_425_0_sva <= sigmoid_table_425_0_sva_dfm_1;
      sigmoid_table_425_4_sva <= sigmoid_table_425_4_sva_dfm_1;
      sigmoid_table_422_0_sva <= sigmoid_table_422_0_sva_dfm_1;
      sigmoid_table_422_3_sva <= sigmoid_table_422_3_sva_dfm_1;
      sigmoid_table_420_2_sva <= sigmoid_table_420_2_sva_dfm_1;
      sigmoid_table_419_1_sva <= sigmoid_table_419_1_sva_dfm_1;
      sigmoid_table_418_7_sva <= sigmoid_table_418_7_sva_dfm_1;
      sigmoid_table_417_0_sva <= sigmoid_table_417_0_sva_dfm_1;
      sigmoid_table_417_7_sva <= sigmoid_table_417_7_sva_dfm_1;
      sigmoid_table_416_1_sva <= sigmoid_table_416_1_sva_dfm_1;
      sigmoid_table_416_7_sva <= sigmoid_table_416_7_sva_dfm_1;
      sigmoid_table_415_7_sva <= sigmoid_table_415_7_sva_dfm_1;
      sigmoid_table_414_7_sva <= sigmoid_table_414_7_sva_dfm_1;
      sigmoid_table_413_7_sva <= sigmoid_table_413_7_sva_dfm_1;
      sigmoid_table_412_0_sva <= sigmoid_table_412_0_sva_dfm_1;
      sigmoid_table_412_7_sva <= sigmoid_table_412_7_sva_dfm_1;
      sigmoid_table_411_5_sva <= sigmoid_table_411_5_sva_dfm_1;
      sigmoid_table_411_7_sva <= sigmoid_table_411_7_sva_dfm_1;
      sigmoid_table_410_5_sva <= sigmoid_table_410_5_sva_dfm_1;
      sigmoid_table_410_7_sva <= sigmoid_table_410_7_sva_dfm_1;
      sigmoid_table_409_1_sva <= sigmoid_table_409_1_sva_dfm_1;
      sigmoid_table_409_3_sva <= sigmoid_table_409_3_sva_dfm_1;
      sigmoid_table_409_5_sva <= sigmoid_table_409_5_sva_dfm_1;
      sigmoid_table_409_7_sva <= sigmoid_table_409_7_sva_dfm_1;
      sigmoid_table_408_3_sva <= sigmoid_table_408_3_sva_dfm_1;
      sigmoid_table_408_5_sva <= sigmoid_table_408_5_sva_dfm_1;
      sigmoid_table_408_7_sva <= sigmoid_table_408_7_sva_dfm_1;
      sigmoid_table_407_5_sva <= sigmoid_table_407_5_sva_dfm_1;
      sigmoid_table_407_7_sva <= sigmoid_table_407_7_sva_dfm_1;
      sigmoid_table_406_2_sva <= sigmoid_table_406_2_sva_dfm_1;
      sigmoid_table_406_5_sva <= sigmoid_table_406_5_sva_dfm_1;
      sigmoid_table_406_7_sva <= sigmoid_table_406_7_sva_dfm_1;
      sigmoid_table_405_0_sva <= sigmoid_table_405_0_sva_dfm_1;
      sigmoid_table_405_5_sva <= sigmoid_table_405_5_sva_dfm_1;
      sigmoid_table_405_7_sva <= sigmoid_table_405_7_sva_dfm_1;
      sigmoid_table_404_7_sva <= sigmoid_table_404_7_sva_dfm_1;
      sigmoid_table_403_0_sva <= sigmoid_table_403_0_sva_dfm_1;
      sigmoid_table_403_7_sva <= sigmoid_table_403_7_sva_dfm_1;
      sigmoid_table_402_7_sva <= sigmoid_table_402_7_sva_dfm_1;
      sigmoid_table_401_0_sva <= sigmoid_table_401_0_sva_dfm_1;
      sigmoid_table_401_7_sva <= sigmoid_table_401_7_sva_dfm_1;
      sigmoid_table_400_4_sva <= sigmoid_table_400_4_sva_dfm_1;
      sigmoid_table_400_7_sva <= sigmoid_table_400_7_sva_dfm_1;
      sigmoid_table_399_0_sva <= sigmoid_table_399_0_sva_dfm_1;
      sigmoid_table_399_2_sva <= sigmoid_table_399_2_sva_dfm_1;
      sigmoid_table_399_4_sva <= sigmoid_table_399_4_sva_dfm_1;
      sigmoid_table_399_7_sva <= sigmoid_table_399_7_sva_dfm_1;
      sigmoid_table_398_4_sva <= sigmoid_table_398_4_sva_dfm_1;
      sigmoid_table_398_7_sva <= sigmoid_table_398_7_sva_dfm_1;
      sigmoid_table_397_0_sva <= sigmoid_table_397_0_sva_dfm_1;
      sigmoid_table_397_4_sva <= sigmoid_table_397_4_sva_dfm_1;
      sigmoid_table_397_7_sva <= sigmoid_table_397_7_sva_dfm_1;
      sigmoid_table_396_7_sva <= sigmoid_table_396_7_sva_dfm_1;
      sigmoid_table_395_0_sva <= sigmoid_table_395_0_sva_dfm_1;
      sigmoid_table_395_7_sva <= sigmoid_table_395_7_sva_dfm_1;
      sigmoid_table_394_3_sva <= sigmoid_table_394_3_sva_dfm_1;
      sigmoid_table_394_7_sva <= sigmoid_table_394_7_sva_dfm_1;
      sigmoid_table_393_1_sva <= sigmoid_table_393_1_sva_dfm_1;
      sigmoid_table_393_3_sva <= sigmoid_table_393_3_sva_dfm_1;
      sigmoid_table_393_7_sva <= sigmoid_table_393_7_sva_dfm_1;
      sigmoid_table_392_3_sva <= sigmoid_table_392_3_sva_dfm_1;
      sigmoid_table_392_7_sva <= sigmoid_table_392_7_sva_dfm_1;
      sigmoid_table_391_7_sva <= sigmoid_table_391_7_sva_dfm_1;
      sigmoid_table_390_2_sva <= sigmoid_table_390_2_sva_dfm_1;
      sigmoid_table_390_7_sva <= sigmoid_table_390_7_sva_dfm_1;
      sigmoid_table_389_1_sva <= sigmoid_table_389_1_sva_dfm_1;
      sigmoid_table_389_7_sva <= sigmoid_table_389_7_sva_dfm_1;
      sigmoid_table_388_7_sva <= sigmoid_table_388_7_sva_dfm_1;
      sigmoid_table_386_0_sva <= sigmoid_table_386_0_sva_dfm_1;
      sigmoid_table_384_1_sva <= sigmoid_table_384_1_sva_dfm_1;
      sigmoid_table_381_0_sva <= sigmoid_table_381_0_sva_dfm_1;
      sigmoid_table_381_2_sva <= sigmoid_table_381_2_sva_dfm_1;
      sigmoid_table_379_0_sva <= sigmoid_table_379_0_sva_dfm_1;
      sigmoid_table_376_0_sva <= sigmoid_table_376_0_sva_dfm_1;
      sigmoid_table_375_3_sva <= sigmoid_table_375_3_sva_dfm_1;
      sigmoid_table_374_1_sva <= sigmoid_table_374_1_sva_dfm_1;
      sigmoid_table_374_3_sva <= sigmoid_table_374_3_sva_dfm_1;
      sigmoid_table_373_3_sva <= sigmoid_table_373_3_sva_dfm_1;
      sigmoid_table_371_0_sva <= sigmoid_table_371_0_sva_dfm_1;
      sigmoid_table_371_2_sva <= sigmoid_table_371_2_sva_dfm_1;
      sigmoid_table_370_2_sva <= sigmoid_table_370_2_sva_dfm_1;
      sigmoid_table_368_0_sva <= sigmoid_table_368_0_sva_dfm_1;
      sigmoid_table_366_6_sva <= sigmoid_table_366_6_sva_dfm_1;
      sigmoid_table_365_0_sva <= sigmoid_table_365_0_sva_dfm_1;
      sigmoid_table_365_6_sva <= sigmoid_table_365_6_sva_dfm_1;
      sigmoid_table_364_6_sva <= sigmoid_table_364_6_sva_dfm_1;
      sigmoid_table_363_1_sva <= sigmoid_table_363_1_sva_dfm_1;
      sigmoid_table_363_6_sva <= sigmoid_table_363_6_sva_dfm_1;
      sigmoid_table_362_0_sva <= sigmoid_table_362_0_sva_dfm_1;
      sigmoid_table_362_6_sva <= sigmoid_table_362_6_sva_dfm_1;
      sigmoid_table_361_6_sva <= sigmoid_table_361_6_sva_dfm_1;
      sigmoid_table_360_4_sva <= sigmoid_table_360_4_sva_dfm_1;
      sigmoid_table_360_6_sva <= sigmoid_table_360_6_sva_dfm_1;
      sigmoid_table_359_0_sva <= sigmoid_table_359_0_sva_dfm_1;
      sigmoid_table_359_2_sva <= sigmoid_table_359_2_sva_dfm_1;
      sigmoid_table_359_4_sva <= sigmoid_table_359_4_sva_dfm_1;
      sigmoid_table_359_6_sva <= sigmoid_table_359_6_sva_dfm_1;
      sigmoid_table_358_2_sva <= sigmoid_table_358_2_sva_dfm_1;
      sigmoid_table_358_4_sva <= sigmoid_table_358_4_sva_dfm_1;
      sigmoid_table_358_6_sva <= sigmoid_table_358_6_sva_dfm_1;
      sigmoid_table_357_4_sva <= sigmoid_table_357_4_sva_dfm_1;
      sigmoid_table_357_6_sva <= sigmoid_table_357_6_sva_dfm_1;
      sigmoid_table_356_1_sva <= sigmoid_table_356_1_sva_dfm_1;
      sigmoid_table_356_4_sva <= sigmoid_table_356_4_sva_dfm_1;
      sigmoid_table_356_6_sva <= sigmoid_table_356_6_sva_dfm_1;
      sigmoid_table_355_0_sva <= sigmoid_table_355_0_sva_dfm_1;
      sigmoid_table_355_4_sva <= sigmoid_table_355_4_sva_dfm_1;
      sigmoid_table_355_6_sva <= sigmoid_table_355_6_sva_dfm_1;
      sigmoid_table_354_6_sva <= sigmoid_table_354_6_sva_dfm_1;
      sigmoid_table_353_6_sva <= sigmoid_table_353_6_sva_dfm_1;
      sigmoid_table_352_0_sva <= sigmoid_table_352_0_sva_dfm_1;
      sigmoid_table_352_6_sva <= sigmoid_table_352_6_sva_dfm_1;
      sigmoid_table_351_6_sva <= sigmoid_table_351_6_sva_dfm_1;
      sigmoid_table_350_3_sva <= sigmoid_table_350_3_sva_dfm_1;
      sigmoid_table_350_6_sva <= sigmoid_table_350_6_sva_dfm_1;
      sigmoid_table_349_1_sva <= sigmoid_table_349_1_sva_dfm_1;
      sigmoid_table_349_3_sva <= sigmoid_table_349_3_sva_dfm_1;
      sigmoid_table_349_6_sva <= sigmoid_table_349_6_sva_dfm_1;
      sigmoid_table_348_0_sva <= sigmoid_table_348_0_sva_dfm_1;
      sigmoid_table_348_3_sva <= sigmoid_table_348_3_sva_dfm_1;
      sigmoid_table_348_6_sva <= sigmoid_table_348_6_sva_dfm_1;
      sigmoid_table_347_3_sva <= sigmoid_table_347_3_sva_dfm_1;
      sigmoid_table_347_6_sva <= sigmoid_table_347_6_sva_dfm_1;
      sigmoid_table_346_6_sva <= sigmoid_table_346_6_sva_dfm_1;
      sigmoid_table_345_6_sva <= sigmoid_table_345_6_sva_dfm_1;
      sigmoid_table_344_0_sva <= sigmoid_table_344_0_sva_dfm_1;
      sigmoid_table_344_2_sva <= sigmoid_table_344_2_sva_dfm_1;
      sigmoid_table_344_6_sva <= sigmoid_table_344_6_sva_dfm_1;
      sigmoid_table_343_2_sva <= sigmoid_table_343_2_sva_dfm_1;
      sigmoid_table_343_6_sva <= sigmoid_table_343_6_sva_dfm_1;
      sigmoid_table_342_6_sva <= sigmoid_table_342_6_sva_dfm_1;
      sigmoid_table_341_1_sva <= sigmoid_table_341_1_sva_dfm_1;
      sigmoid_table_341_6_sva <= sigmoid_table_341_6_sva_dfm_1;
      sigmoid_table_340_0_sva <= sigmoid_table_340_0_sva_dfm_1;
      sigmoid_table_340_6_sva <= sigmoid_table_340_6_sva_dfm_1;
      sigmoid_table_339_6_sva <= sigmoid_table_339_6_sva_dfm_1;
      sigmoid_table_336_0_sva <= sigmoid_table_336_0_sva_dfm_1;
      sigmoid_table_333_1_sva <= sigmoid_table_333_1_sva_dfm_1;
      sigmoid_table_332_1_sva <= sigmoid_table_332_1_sva_dfm_1;
      sigmoid_table_331_0_sva <= sigmoid_table_331_0_sva_dfm_1;
      sigmoid_table_327_0_sva <= sigmoid_table_327_0_sva_dfm_1;
      sigmoid_table_327_2_sva <= sigmoid_table_327_2_sva_dfm_1;
      sigmoid_table_326_0_sva <= sigmoid_table_326_0_sva_dfm_1;
      sigmoid_table_326_2_sva <= sigmoid_table_326_2_sva_dfm_1;
      sigmoid_table_325_2_sva <= sigmoid_table_325_2_sva_dfm_1;
      sigmoid_table_323_1_sva <= sigmoid_table_323_1_sva_dfm_1;
      sigmoid_table_322_1_sva <= sigmoid_table_322_1_sva_dfm_1;
      sigmoid_table_321_0_sva <= sigmoid_table_321_0_sva_dfm_1;
      sigmoid_table_319_5_sva <= sigmoid_table_319_5_sva_dfm_1;
      sigmoid_table_318_5_sva <= sigmoid_table_318_5_sva_dfm_1;
      sigmoid_table_317_5_sva <= sigmoid_table_317_5_sva_dfm_1;
      sigmoid_table_316_0_sva <= sigmoid_table_316_0_sva_dfm_1;
      sigmoid_table_316_5_sva <= sigmoid_table_316_5_sva_dfm_1;
      sigmoid_table_315_0_sva <= sigmoid_table_315_0_sva_dfm_1;
      sigmoid_table_315_5_sva <= sigmoid_table_315_5_sva_dfm_1;
      sigmoid_table_314_5_sva <= sigmoid_table_314_5_sva_dfm_1;
      sigmoid_table_313_3_sva <= sigmoid_table_313_3_sva_dfm_1;
      sigmoid_table_313_5_sva <= sigmoid_table_313_5_sva_dfm_1;
      sigmoid_table_312_3_sva <= sigmoid_table_312_3_sva_dfm_1;
      sigmoid_table_312_5_sva <= sigmoid_table_312_5_sva_dfm_1;
      sigmoid_table_311_1_sva <= sigmoid_table_311_1_sva_dfm_1;
      sigmoid_table_311_3_sva <= sigmoid_table_311_3_sva_dfm_1;
      sigmoid_table_311_5_sva <= sigmoid_table_311_5_sva_dfm_1;
      sigmoid_table_310_0_sva <= sigmoid_table_310_0_sva_dfm_1;
      sigmoid_table_310_3_sva <= sigmoid_table_310_3_sva_dfm_1;
      sigmoid_table_310_5_sva <= sigmoid_table_310_5_sva_dfm_1;
      sigmoid_table_309_0_sva <= sigmoid_table_309_0_sva_dfm_1;
      sigmoid_table_309_3_sva <= sigmoid_table_309_3_sva_dfm_1;
      sigmoid_table_309_5_sva <= sigmoid_table_309_5_sva_dfm_1;
      sigmoid_table_308_3_sva <= sigmoid_table_308_3_sva_dfm_1;
      sigmoid_table_308_5_sva <= sigmoid_table_308_5_sva_dfm_1;
      sigmoid_table_307_5_sva <= sigmoid_table_307_5_sva_dfm_1;
      sigmoid_table_306_5_sva <= sigmoid_table_306_5_sva_dfm_1;
      sigmoid_table_305_5_sva <= sigmoid_table_305_5_sva_dfm_1;
      sigmoid_table_304_5_sva <= sigmoid_table_304_5_sva_dfm_1;
      sigmoid_table_303_0_sva <= sigmoid_table_303_0_sva_dfm_1;
      sigmoid_table_303_2_sva <= sigmoid_table_303_2_sva_dfm_1;
      sigmoid_table_303_5_sva <= sigmoid_table_303_5_sva_dfm_1;
      sigmoid_table_302_0_sva <= sigmoid_table_302_0_sva_dfm_1;
      sigmoid_table_302_2_sva <= sigmoid_table_302_2_sva_dfm_1;
      sigmoid_table_302_5_sva <= sigmoid_table_302_5_sva_dfm_1;
      sigmoid_table_301_2_sva <= sigmoid_table_301_2_sva_dfm_1;
      sigmoid_table_301_5_sva <= sigmoid_table_301_5_sva_dfm_1;
      sigmoid_table_300_5_sva <= sigmoid_table_300_5_sva_dfm_1;
      sigmoid_table_299_5_sva <= sigmoid_table_299_5_sva_dfm_1;
      sigmoid_table_298_1_sva <= sigmoid_table_298_1_sva_dfm_1;
      sigmoid_table_298_5_sva <= sigmoid_table_298_5_sva_dfm_1;
      sigmoid_table_297_1_sva <= sigmoid_table_297_1_sva_dfm_1;
      sigmoid_table_297_5_sva <= sigmoid_table_297_5_sva_dfm_1;
      sigmoid_table_296_0_sva <= sigmoid_table_296_0_sva_dfm_1;
      sigmoid_table_296_5_sva <= sigmoid_table_296_5_sva_dfm_1;
      sigmoid_table_295_0_sva <= sigmoid_table_295_0_sva_dfm_1;
      sigmoid_table_295_5_sva <= sigmoid_table_295_5_sva_dfm_1;
      sigmoid_table_294_5_sva <= sigmoid_table_294_5_sva_dfm_1;
      sigmoid_table_293_5_sva <= sigmoid_table_293_5_sva_dfm_1;
      sigmoid_table_287_0_sva <= sigmoid_table_287_0_sva_dfm_1;
      sigmoid_table_286_0_sva <= sigmoid_table_286_0_sva_dfm_1;
      sigmoid_table_281_1_sva <= sigmoid_table_281_1_sva_dfm_1;
      sigmoid_table_280_1_sva <= sigmoid_table_280_1_sva_dfm_1;
      sigmoid_table_279_1_sva <= sigmoid_table_279_1_sva_dfm_1;
      sigmoid_table_278_0_sva <= sigmoid_table_278_0_sva_dfm_1;
      sigmoid_table_277_0_sva <= sigmoid_table_277_0_sva_dfm_1;
      sigmoid_table_276_0_sva <= sigmoid_table_276_0_sva_dfm_1;
      sigmoid_table_273_4_sva <= sigmoid_table_273_4_sva_dfm_1;
      sigmoid_table_272_4_sva <= sigmoid_table_272_4_sva_dfm_1;
      sigmoid_table_271_4_sva <= sigmoid_table_271_4_sva_dfm_1;
      sigmoid_table_270_4_sva <= sigmoid_table_270_4_sva_dfm_1;
      sigmoid_table_269_4_sva <= sigmoid_table_269_4_sva_dfm_1;
      sigmoid_table_268_4_sva <= sigmoid_table_268_4_sva_dfm_1;
      sigmoid_table_267_0_sva <= sigmoid_table_267_0_sva_dfm_1;
      sigmoid_table_267_2_sva <= sigmoid_table_267_2_sva_dfm_1;
      sigmoid_table_267_4_sva <= sigmoid_table_267_4_sva_dfm_1;
      sigmoid_table_266_0_sva <= sigmoid_table_266_0_sva_dfm_1;
      sigmoid_table_266_2_sva <= sigmoid_table_266_2_sva_dfm_1;
      sigmoid_table_266_4_sva <= sigmoid_table_266_4_sva_dfm_1;
      sigmoid_table_265_0_sva <= sigmoid_table_265_0_sva_dfm_1;
      sigmoid_table_265_2_sva <= sigmoid_table_265_2_sva_dfm_1;
      sigmoid_table_265_4_sva <= sigmoid_table_265_4_sva_dfm_1;
      sigmoid_table_264_2_sva <= sigmoid_table_264_2_sva_dfm_1;
      sigmoid_table_264_4_sva <= sigmoid_table_264_4_sva_dfm_1;
      sigmoid_table_263_2_sva <= sigmoid_table_263_2_sva_dfm_1;
      sigmoid_table_263_4_sva <= sigmoid_table_263_4_sva_dfm_1;
      sigmoid_table_262_2_sva <= sigmoid_table_262_2_sva_dfm_1;
      sigmoid_table_262_4_sva <= sigmoid_table_262_4_sva_dfm_1;
      sigmoid_table_261_4_sva <= sigmoid_table_261_4_sva_dfm_1;
      sigmoid_table_260_4_sva <= sigmoid_table_260_4_sva_dfm_1;
      sigmoid_table_259_4_sva <= sigmoid_table_259_4_sva_dfm_1;
      sigmoid_table_258_1_sva <= sigmoid_table_258_1_sva_dfm_1;
      sigmoid_table_258_4_sva <= sigmoid_table_258_4_sva_dfm_1;
      sigmoid_table_257_1_sva <= sigmoid_table_257_1_sva_dfm_1;
      sigmoid_table_257_4_sva <= sigmoid_table_257_4_sva_dfm_1;
      sigmoid_table_256_1_sva <= sigmoid_table_256_1_sva_dfm_1;
      sigmoid_table_256_4_sva <= sigmoid_table_256_4_sva_dfm_1;
      sigmoid_table_255_1_sva <= sigmoid_table_255_1_sva_dfm_1;
      sigmoid_table_255_4_sva <= sigmoid_table_255_4_sva_dfm_1;
      sigmoid_table_254_0_sva <= sigmoid_table_254_0_sva_dfm_1;
      sigmoid_table_254_4_sva <= sigmoid_table_254_4_sva_dfm_1;
      sigmoid_table_253_0_sva <= sigmoid_table_253_0_sva_dfm_1;
      sigmoid_table_253_4_sva <= sigmoid_table_253_4_sva_dfm_1;
      sigmoid_table_252_0_sva <= sigmoid_table_252_0_sva_dfm_1;
      sigmoid_table_252_4_sva <= sigmoid_table_252_4_sva_dfm_1;
      sigmoid_table_251_0_sva <= sigmoid_table_251_0_sva_dfm_1;
      sigmoid_table_251_4_sva <= sigmoid_table_251_4_sva_dfm_1;
      sigmoid_table_250_4_sva <= sigmoid_table_250_4_sva_dfm_1;
      sigmoid_table_249_4_sva <= sigmoid_table_249_4_sva_dfm_1;
      sigmoid_table_248_4_sva <= sigmoid_table_248_4_sva_dfm_1;
      sigmoid_table_247_4_sva <= sigmoid_table_247_4_sva_dfm_1;
      sigmoid_table_238_0_sva <= sigmoid_table_238_0_sva_dfm_1;
      sigmoid_table_237_0_sva <= sigmoid_table_237_0_sva_dfm_1;
      sigmoid_table_236_0_sva <= sigmoid_table_236_0_sva_dfm_1;
      sigmoid_table_235_0_sva <= sigmoid_table_235_0_sva_dfm_1;
      sigmoid_table_234_0_sva <= sigmoid_table_234_0_sva_dfm_1;
      sigmoid_table_228_3_sva <= sigmoid_table_228_3_sva_dfm_1;
      sigmoid_table_227_3_sva <= sigmoid_table_227_3_sva_dfm_1;
      sigmoid_table_226_3_sva <= sigmoid_table_226_3_sva_dfm_1;
      sigmoid_table_225_3_sva <= sigmoid_table_225_3_sva_dfm_1;
      sigmoid_table_224_3_sva <= sigmoid_table_224_3_sva_dfm_1;
      sigmoid_table_223_3_sva <= sigmoid_table_223_3_sva_dfm_1;
      sigmoid_table_222_1_sva <= sigmoid_table_222_1_sva_dfm_1;
      sigmoid_table_222_3_sva <= sigmoid_table_222_3_sva_dfm_1;
      sigmoid_table_221_1_sva <= sigmoid_table_221_1_sva_dfm_1;
      sigmoid_table_221_3_sva <= sigmoid_table_221_3_sva_dfm_1;
      sigmoid_table_220_1_sva <= sigmoid_table_220_1_sva_dfm_1;
      sigmoid_table_220_3_sva <= sigmoid_table_220_3_sva_dfm_1;
      sigmoid_table_219_1_sva <= sigmoid_table_219_1_sva_dfm_1;
      sigmoid_table_219_3_sva <= sigmoid_table_219_3_sva_dfm_1;
      sigmoid_table_218_1_sva <= sigmoid_table_218_1_sva_dfm_1;
      sigmoid_table_218_3_sva <= sigmoid_table_218_3_sva_dfm_1;
      sigmoid_table_217_1_sva <= sigmoid_table_217_1_sva_dfm_1;
      sigmoid_table_217_3_sva <= sigmoid_table_217_3_sva_dfm_1;
      sigmoid_table_216_0_sva <= sigmoid_table_216_0_sva_dfm_1;
      sigmoid_table_216_3_sva <= sigmoid_table_216_3_sva_dfm_1;
      sigmoid_table_215_0_sva <= sigmoid_table_215_0_sva_dfm_1;
      sigmoid_table_215_3_sva <= sigmoid_table_215_3_sva_dfm_1;
      sigmoid_table_214_0_sva <= sigmoid_table_214_0_sva_dfm_1;
      sigmoid_table_214_3_sva <= sigmoid_table_214_3_sva_dfm_1;
      sigmoid_table_213_0_sva <= sigmoid_table_213_0_sva_dfm_1;
      sigmoid_table_213_3_sva <= sigmoid_table_213_3_sva_dfm_1;
      sigmoid_table_212_0_sva <= sigmoid_table_212_0_sva_dfm_1;
      sigmoid_table_212_3_sva <= sigmoid_table_212_3_sva_dfm_1;
      sigmoid_table_211_0_sva <= sigmoid_table_211_0_sva_dfm_1;
      sigmoid_table_211_3_sva <= sigmoid_table_211_3_sva_dfm_1;
      sigmoid_table_210_0_sva <= sigmoid_table_210_0_sva_dfm_1;
      sigmoid_table_210_3_sva <= sigmoid_table_210_3_sva_dfm_1;
      sigmoid_table_209_3_sva <= sigmoid_table_209_3_sva_dfm_1;
      sigmoid_table_208_3_sva <= sigmoid_table_208_3_sva_dfm_1;
      sigmoid_table_207_3_sva <= sigmoid_table_207_3_sva_dfm_1;
      sigmoid_table_206_3_sva <= sigmoid_table_206_3_sva_dfm_1;
      sigmoid_table_205_3_sva <= sigmoid_table_205_3_sva_dfm_1;
      sigmoid_table_204_3_sva <= sigmoid_table_204_3_sva_dfm_1;
      sigmoid_table_203_3_sva <= sigmoid_table_203_3_sva_dfm_1;
      sigmoid_table_202_3_sva <= sigmoid_table_202_3_sva_dfm_1;
      sigmoid_table_183_0_sva <= sigmoid_table_183_0_sva_dfm_1;
      sigmoid_table_183_2_sva <= sigmoid_table_183_2_sva_dfm_1;
      sigmoid_table_182_0_sva <= sigmoid_table_182_0_sva_dfm_1;
      sigmoid_table_182_2_sva <= sigmoid_table_182_2_sva_dfm_1;
      sigmoid_table_181_0_sva <= sigmoid_table_181_0_sva_dfm_1;
      sigmoid_table_181_2_sva <= sigmoid_table_181_2_sva_dfm_1;
      sigmoid_table_180_0_sva <= sigmoid_table_180_0_sva_dfm_1;
      sigmoid_table_180_2_sva <= sigmoid_table_180_2_sva_dfm_1;
      sigmoid_table_179_0_sva <= sigmoid_table_179_0_sva_dfm_1;
      sigmoid_table_179_2_sva <= sigmoid_table_179_2_sva_dfm_1;
      sigmoid_table_178_0_sva <= sigmoid_table_178_0_sva_dfm_1;
      sigmoid_table_178_2_sva <= sigmoid_table_178_2_sva_dfm_1;
      sigmoid_table_177_0_sva <= sigmoid_table_177_0_sva_dfm_1;
      sigmoid_table_177_2_sva <= sigmoid_table_177_2_sva_dfm_1;
      sigmoid_table_176_0_sva <= sigmoid_table_176_0_sva_dfm_1;
      sigmoid_table_176_2_sva <= sigmoid_table_176_2_sva_dfm_1;
      sigmoid_table_175_0_sva <= sigmoid_table_175_0_sva_dfm_1;
      sigmoid_table_175_2_sva <= sigmoid_table_175_2_sva_dfm_1;
      sigmoid_table_174_0_sva <= sigmoid_table_174_0_sva_dfm_1;
      sigmoid_table_174_2_sva <= sigmoid_table_174_2_sva_dfm_1;
      sigmoid_table_173_0_sva <= sigmoid_table_173_0_sva_dfm_1;
      sigmoid_table_173_2_sva <= sigmoid_table_173_2_sva_dfm_1;
      sigmoid_table_172_0_sva <= sigmoid_table_172_0_sva_dfm_1;
      sigmoid_table_172_2_sva <= sigmoid_table_172_2_sva_dfm_1;
      sigmoid_table_171_2_sva <= sigmoid_table_171_2_sva_dfm_1;
      sigmoid_table_170_2_sva <= sigmoid_table_170_2_sva_dfm_1;
      sigmoid_table_169_2_sva <= sigmoid_table_169_2_sva_dfm_1;
      sigmoid_table_168_2_sva <= sigmoid_table_168_2_sva_dfm_1;
      sigmoid_table_167_2_sva <= sigmoid_table_167_2_sva_dfm_1;
      sigmoid_table_166_2_sva <= sigmoid_table_166_2_sva_dfm_1;
      sigmoid_table_165_2_sva <= sigmoid_table_165_2_sva_dfm_1;
      sigmoid_table_164_2_sva <= sigmoid_table_164_2_sva_dfm_1;
      sigmoid_table_163_2_sva <= sigmoid_table_163_2_sva_dfm_1;
      sigmoid_table_162_2_sva <= sigmoid_table_162_2_sva_dfm_1;
      sigmoid_table_161_2_sva <= sigmoid_table_161_2_sva_dfm_1;
      sigmoid_table_160_2_sva <= sigmoid_table_160_2_sva_dfm_1;
      sigmoid_table_159_2_sva <= sigmoid_table_159_2_sva_dfm_1;
      sigmoid_table_158_2_sva <= sigmoid_table_158_2_sva_dfm_1;
      sigmoid_table_138_1_sva <= sigmoid_table_138_1_sva_dfm_1;
      sigmoid_table_137_1_sva <= sigmoid_table_137_1_sva_dfm_1;
      sigmoid_table_136_1_sva <= sigmoid_table_136_1_sva_dfm_1;
      sigmoid_table_135_1_sva <= sigmoid_table_135_1_sva_dfm_1;
      sigmoid_table_134_1_sva <= sigmoid_table_134_1_sva_dfm_1;
      sigmoid_table_133_1_sva <= sigmoid_table_133_1_sva_dfm_1;
      sigmoid_table_132_1_sva <= sigmoid_table_132_1_sva_dfm_1;
      sigmoid_table_131_1_sva <= sigmoid_table_131_1_sva_dfm_1;
      sigmoid_table_130_1_sva <= sigmoid_table_130_1_sva_dfm_1;
      sigmoid_table_129_1_sva <= sigmoid_table_129_1_sva_dfm_1;
      sigmoid_table_128_1_sva <= sigmoid_table_128_1_sva_dfm_1;
      sigmoid_table_127_1_sva <= sigmoid_table_127_1_sva_dfm_1;
      sigmoid_table_126_1_sva <= sigmoid_table_126_1_sva_dfm_1;
      sigmoid_table_125_1_sva <= sigmoid_table_125_1_sva_dfm_1;
      sigmoid_table_124_1_sva <= sigmoid_table_124_1_sva_dfm_1;
      sigmoid_table_123_1_sva <= sigmoid_table_123_1_sva_dfm_1;
      sigmoid_table_122_1_sva <= sigmoid_table_122_1_sva_dfm_1;
      sigmoid_table_121_1_sva <= sigmoid_table_121_1_sva_dfm_1;
      sigmoid_table_120_1_sva <= sigmoid_table_120_1_sva_dfm_1;
      sigmoid_table_119_1_sva <= sigmoid_table_119_1_sva_dfm_1;
      sigmoid_table_118_1_sva <= sigmoid_table_118_1_sva_dfm_1;
      sigmoid_table_117_1_sva <= sigmoid_table_117_1_sva_dfm_1;
      sigmoid_table_116_1_sva <= sigmoid_table_116_1_sva_dfm_1;
      sigmoid_table_115_1_sva <= sigmoid_table_115_1_sva_dfm_1;
      sigmoid_table_114_1_sva <= sigmoid_table_114_1_sva_dfm_1;
      sigmoid_table_113_1_sva <= sigmoid_table_113_1_sva_dfm_1;
      sigmoid_table_112_0_sva <= sigmoid_table_112_0_sva_dfm_1;
      sigmoid_table_111_0_sva <= sigmoid_table_111_0_sva_dfm_1;
      sigmoid_table_110_0_sva <= sigmoid_table_110_0_sva_dfm_1;
      sigmoid_table_109_0_sva <= sigmoid_table_109_0_sva_dfm_1;
      sigmoid_table_108_0_sva <= sigmoid_table_108_0_sva_dfm_1;
      sigmoid_table_107_0_sva <= sigmoid_table_107_0_sva_dfm_1;
      sigmoid_table_106_0_sva <= sigmoid_table_106_0_sva_dfm_1;
      sigmoid_table_105_0_sva <= sigmoid_table_105_0_sva_dfm_1;
      sigmoid_table_104_0_sva <= sigmoid_table_104_0_sva_dfm_1;
      sigmoid_table_103_0_sva <= sigmoid_table_103_0_sva_dfm_1;
      sigmoid_table_102_0_sva <= sigmoid_table_102_0_sva_dfm_1;
      sigmoid_table_101_0_sva <= sigmoid_table_101_0_sva_dfm_1;
      sigmoid_table_100_0_sva <= sigmoid_table_100_0_sva_dfm_1;
      sigmoid_table_99_0_sva <= sigmoid_table_99_0_sva_dfm_1;
      sigmoid_table_98_0_sva <= sigmoid_table_98_0_sva_dfm_1;
      sigmoid_table_97_0_sva <= sigmoid_table_97_0_sva_dfm_1;
      sigmoid_table_96_0_sva <= sigmoid_table_96_0_sva_dfm_1;
      sigmoid_table_95_0_sva <= sigmoid_table_95_0_sva_dfm_1;
      sigmoid_table_94_0_sva <= sigmoid_table_94_0_sva_dfm_1;
      sigmoid_table_93_0_sva <= sigmoid_table_93_0_sva_dfm_1;
      sigmoid_table_92_0_sva <= sigmoid_table_92_0_sva_dfm_1;
      sigmoid_table_91_0_sva <= sigmoid_table_91_0_sva_dfm_1;
      sigmoid_table_90_0_sva <= sigmoid_table_90_0_sva_dfm_1;
      sigmoid_table_89_0_sva <= sigmoid_table_89_0_sva_dfm_1;
      sigmoid_table_88_0_sva <= sigmoid_table_88_0_sva_dfm_1;
      sigmoid_table_87_0_sva <= sigmoid_table_87_0_sva_dfm_1;
      sigmoid_table_86_0_sva <= sigmoid_table_86_0_sva_dfm_1;
      sigmoid_table_85_0_sva <= sigmoid_table_85_0_sva_dfm_1;
      sigmoid_table_84_0_sva <= sigmoid_table_84_0_sva_dfm_1;
      sigmoid_table_83_0_sva <= sigmoid_table_83_0_sva_dfm_1;
      sigmoid_table_82_0_sva <= sigmoid_table_82_0_sva_dfm_1;
      sigmoid_table_81_0_sva <= sigmoid_table_81_0_sva_dfm_1;
      sigmoid_table_80_0_sva <= sigmoid_table_80_0_sva_dfm_1;
      sigmoid_table_79_0_sva <= sigmoid_table_79_0_sva_dfm_1;
      sigmoid_table_78_0_sva <= sigmoid_table_78_0_sva_dfm_1;
      sigmoid_table_77_0_sva <= sigmoid_table_77_0_sva_dfm_1;
      sigmoid_table_76_0_sva <= sigmoid_table_76_0_sva_dfm_1;
      sigmoid_table_75_0_sva <= sigmoid_table_75_0_sva_dfm_1;
      sigmoid_table_74_0_sva <= sigmoid_table_74_0_sva_dfm_1;
      sigmoid_table_73_0_sva <= sigmoid_table_73_0_sva_dfm_1;
      sigmoid_table_72_0_sva <= sigmoid_table_72_0_sva_dfm_1;
      sigmoid_table_71_0_sva <= sigmoid_table_71_0_sva_dfm_1;
      sigmoid_table_70_0_sva <= sigmoid_table_70_0_sva_dfm_1;
      sigmoid_table_69_0_sva <= sigmoid_table_69_0_sva_dfm_1;
    end
  end

  function automatic [0:0] MUX_s_1_1024_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] input_2;
    input [0:0] input_3;
    input [0:0] input_4;
    input [0:0] input_5;
    input [0:0] input_6;
    input [0:0] input_7;
    input [0:0] input_8;
    input [0:0] input_9;
    input [0:0] input_10;
    input [0:0] input_11;
    input [0:0] input_12;
    input [0:0] input_13;
    input [0:0] input_14;
    input [0:0] input_15;
    input [0:0] input_16;
    input [0:0] input_17;
    input [0:0] input_18;
    input [0:0] input_19;
    input [0:0] input_20;
    input [0:0] input_21;
    input [0:0] input_22;
    input [0:0] input_23;
    input [0:0] input_24;
    input [0:0] input_25;
    input [0:0] input_26;
    input [0:0] input_27;
    input [0:0] input_28;
    input [0:0] input_29;
    input [0:0] input_30;
    input [0:0] input_31;
    input [0:0] input_32;
    input [0:0] input_33;
    input [0:0] input_34;
    input [0:0] input_35;
    input [0:0] input_36;
    input [0:0] input_37;
    input [0:0] input_38;
    input [0:0] input_39;
    input [0:0] input_40;
    input [0:0] input_41;
    input [0:0] input_42;
    input [0:0] input_43;
    input [0:0] input_44;
    input [0:0] input_45;
    input [0:0] input_46;
    input [0:0] input_47;
    input [0:0] input_48;
    input [0:0] input_49;
    input [0:0] input_50;
    input [0:0] input_51;
    input [0:0] input_52;
    input [0:0] input_53;
    input [0:0] input_54;
    input [0:0] input_55;
    input [0:0] input_56;
    input [0:0] input_57;
    input [0:0] input_58;
    input [0:0] input_59;
    input [0:0] input_60;
    input [0:0] input_61;
    input [0:0] input_62;
    input [0:0] input_63;
    input [0:0] input_64;
    input [0:0] input_65;
    input [0:0] input_66;
    input [0:0] input_67;
    input [0:0] input_68;
    input [0:0] input_69;
    input [0:0] input_70;
    input [0:0] input_71;
    input [0:0] input_72;
    input [0:0] input_73;
    input [0:0] input_74;
    input [0:0] input_75;
    input [0:0] input_76;
    input [0:0] input_77;
    input [0:0] input_78;
    input [0:0] input_79;
    input [0:0] input_80;
    input [0:0] input_81;
    input [0:0] input_82;
    input [0:0] input_83;
    input [0:0] input_84;
    input [0:0] input_85;
    input [0:0] input_86;
    input [0:0] input_87;
    input [0:0] input_88;
    input [0:0] input_89;
    input [0:0] input_90;
    input [0:0] input_91;
    input [0:0] input_92;
    input [0:0] input_93;
    input [0:0] input_94;
    input [0:0] input_95;
    input [0:0] input_96;
    input [0:0] input_97;
    input [0:0] input_98;
    input [0:0] input_99;
    input [0:0] input_100;
    input [0:0] input_101;
    input [0:0] input_102;
    input [0:0] input_103;
    input [0:0] input_104;
    input [0:0] input_105;
    input [0:0] input_106;
    input [0:0] input_107;
    input [0:0] input_108;
    input [0:0] input_109;
    input [0:0] input_110;
    input [0:0] input_111;
    input [0:0] input_112;
    input [0:0] input_113;
    input [0:0] input_114;
    input [0:0] input_115;
    input [0:0] input_116;
    input [0:0] input_117;
    input [0:0] input_118;
    input [0:0] input_119;
    input [0:0] input_120;
    input [0:0] input_121;
    input [0:0] input_122;
    input [0:0] input_123;
    input [0:0] input_124;
    input [0:0] input_125;
    input [0:0] input_126;
    input [0:0] input_127;
    input [0:0] input_128;
    input [0:0] input_129;
    input [0:0] input_130;
    input [0:0] input_131;
    input [0:0] input_132;
    input [0:0] input_133;
    input [0:0] input_134;
    input [0:0] input_135;
    input [0:0] input_136;
    input [0:0] input_137;
    input [0:0] input_138;
    input [0:0] input_139;
    input [0:0] input_140;
    input [0:0] input_141;
    input [0:0] input_142;
    input [0:0] input_143;
    input [0:0] input_144;
    input [0:0] input_145;
    input [0:0] input_146;
    input [0:0] input_147;
    input [0:0] input_148;
    input [0:0] input_149;
    input [0:0] input_150;
    input [0:0] input_151;
    input [0:0] input_152;
    input [0:0] input_153;
    input [0:0] input_154;
    input [0:0] input_155;
    input [0:0] input_156;
    input [0:0] input_157;
    input [0:0] input_158;
    input [0:0] input_159;
    input [0:0] input_160;
    input [0:0] input_161;
    input [0:0] input_162;
    input [0:0] input_163;
    input [0:0] input_164;
    input [0:0] input_165;
    input [0:0] input_166;
    input [0:0] input_167;
    input [0:0] input_168;
    input [0:0] input_169;
    input [0:0] input_170;
    input [0:0] input_171;
    input [0:0] input_172;
    input [0:0] input_173;
    input [0:0] input_174;
    input [0:0] input_175;
    input [0:0] input_176;
    input [0:0] input_177;
    input [0:0] input_178;
    input [0:0] input_179;
    input [0:0] input_180;
    input [0:0] input_181;
    input [0:0] input_182;
    input [0:0] input_183;
    input [0:0] input_184;
    input [0:0] input_185;
    input [0:0] input_186;
    input [0:0] input_187;
    input [0:0] input_188;
    input [0:0] input_189;
    input [0:0] input_190;
    input [0:0] input_191;
    input [0:0] input_192;
    input [0:0] input_193;
    input [0:0] input_194;
    input [0:0] input_195;
    input [0:0] input_196;
    input [0:0] input_197;
    input [0:0] input_198;
    input [0:0] input_199;
    input [0:0] input_200;
    input [0:0] input_201;
    input [0:0] input_202;
    input [0:0] input_203;
    input [0:0] input_204;
    input [0:0] input_205;
    input [0:0] input_206;
    input [0:0] input_207;
    input [0:0] input_208;
    input [0:0] input_209;
    input [0:0] input_210;
    input [0:0] input_211;
    input [0:0] input_212;
    input [0:0] input_213;
    input [0:0] input_214;
    input [0:0] input_215;
    input [0:0] input_216;
    input [0:0] input_217;
    input [0:0] input_218;
    input [0:0] input_219;
    input [0:0] input_220;
    input [0:0] input_221;
    input [0:0] input_222;
    input [0:0] input_223;
    input [0:0] input_224;
    input [0:0] input_225;
    input [0:0] input_226;
    input [0:0] input_227;
    input [0:0] input_228;
    input [0:0] input_229;
    input [0:0] input_230;
    input [0:0] input_231;
    input [0:0] input_232;
    input [0:0] input_233;
    input [0:0] input_234;
    input [0:0] input_235;
    input [0:0] input_236;
    input [0:0] input_237;
    input [0:0] input_238;
    input [0:0] input_239;
    input [0:0] input_240;
    input [0:0] input_241;
    input [0:0] input_242;
    input [0:0] input_243;
    input [0:0] input_244;
    input [0:0] input_245;
    input [0:0] input_246;
    input [0:0] input_247;
    input [0:0] input_248;
    input [0:0] input_249;
    input [0:0] input_250;
    input [0:0] input_251;
    input [0:0] input_252;
    input [0:0] input_253;
    input [0:0] input_254;
    input [0:0] input_255;
    input [0:0] input_256;
    input [0:0] input_257;
    input [0:0] input_258;
    input [0:0] input_259;
    input [0:0] input_260;
    input [0:0] input_261;
    input [0:0] input_262;
    input [0:0] input_263;
    input [0:0] input_264;
    input [0:0] input_265;
    input [0:0] input_266;
    input [0:0] input_267;
    input [0:0] input_268;
    input [0:0] input_269;
    input [0:0] input_270;
    input [0:0] input_271;
    input [0:0] input_272;
    input [0:0] input_273;
    input [0:0] input_274;
    input [0:0] input_275;
    input [0:0] input_276;
    input [0:0] input_277;
    input [0:0] input_278;
    input [0:0] input_279;
    input [0:0] input_280;
    input [0:0] input_281;
    input [0:0] input_282;
    input [0:0] input_283;
    input [0:0] input_284;
    input [0:0] input_285;
    input [0:0] input_286;
    input [0:0] input_287;
    input [0:0] input_288;
    input [0:0] input_289;
    input [0:0] input_290;
    input [0:0] input_291;
    input [0:0] input_292;
    input [0:0] input_293;
    input [0:0] input_294;
    input [0:0] input_295;
    input [0:0] input_296;
    input [0:0] input_297;
    input [0:0] input_298;
    input [0:0] input_299;
    input [0:0] input_300;
    input [0:0] input_301;
    input [0:0] input_302;
    input [0:0] input_303;
    input [0:0] input_304;
    input [0:0] input_305;
    input [0:0] input_306;
    input [0:0] input_307;
    input [0:0] input_308;
    input [0:0] input_309;
    input [0:0] input_310;
    input [0:0] input_311;
    input [0:0] input_312;
    input [0:0] input_313;
    input [0:0] input_314;
    input [0:0] input_315;
    input [0:0] input_316;
    input [0:0] input_317;
    input [0:0] input_318;
    input [0:0] input_319;
    input [0:0] input_320;
    input [0:0] input_321;
    input [0:0] input_322;
    input [0:0] input_323;
    input [0:0] input_324;
    input [0:0] input_325;
    input [0:0] input_326;
    input [0:0] input_327;
    input [0:0] input_328;
    input [0:0] input_329;
    input [0:0] input_330;
    input [0:0] input_331;
    input [0:0] input_332;
    input [0:0] input_333;
    input [0:0] input_334;
    input [0:0] input_335;
    input [0:0] input_336;
    input [0:0] input_337;
    input [0:0] input_338;
    input [0:0] input_339;
    input [0:0] input_340;
    input [0:0] input_341;
    input [0:0] input_342;
    input [0:0] input_343;
    input [0:0] input_344;
    input [0:0] input_345;
    input [0:0] input_346;
    input [0:0] input_347;
    input [0:0] input_348;
    input [0:0] input_349;
    input [0:0] input_350;
    input [0:0] input_351;
    input [0:0] input_352;
    input [0:0] input_353;
    input [0:0] input_354;
    input [0:0] input_355;
    input [0:0] input_356;
    input [0:0] input_357;
    input [0:0] input_358;
    input [0:0] input_359;
    input [0:0] input_360;
    input [0:0] input_361;
    input [0:0] input_362;
    input [0:0] input_363;
    input [0:0] input_364;
    input [0:0] input_365;
    input [0:0] input_366;
    input [0:0] input_367;
    input [0:0] input_368;
    input [0:0] input_369;
    input [0:0] input_370;
    input [0:0] input_371;
    input [0:0] input_372;
    input [0:0] input_373;
    input [0:0] input_374;
    input [0:0] input_375;
    input [0:0] input_376;
    input [0:0] input_377;
    input [0:0] input_378;
    input [0:0] input_379;
    input [0:0] input_380;
    input [0:0] input_381;
    input [0:0] input_382;
    input [0:0] input_383;
    input [0:0] input_384;
    input [0:0] input_385;
    input [0:0] input_386;
    input [0:0] input_387;
    input [0:0] input_388;
    input [0:0] input_389;
    input [0:0] input_390;
    input [0:0] input_391;
    input [0:0] input_392;
    input [0:0] input_393;
    input [0:0] input_394;
    input [0:0] input_395;
    input [0:0] input_396;
    input [0:0] input_397;
    input [0:0] input_398;
    input [0:0] input_399;
    input [0:0] input_400;
    input [0:0] input_401;
    input [0:0] input_402;
    input [0:0] input_403;
    input [0:0] input_404;
    input [0:0] input_405;
    input [0:0] input_406;
    input [0:0] input_407;
    input [0:0] input_408;
    input [0:0] input_409;
    input [0:0] input_410;
    input [0:0] input_411;
    input [0:0] input_412;
    input [0:0] input_413;
    input [0:0] input_414;
    input [0:0] input_415;
    input [0:0] input_416;
    input [0:0] input_417;
    input [0:0] input_418;
    input [0:0] input_419;
    input [0:0] input_420;
    input [0:0] input_421;
    input [0:0] input_422;
    input [0:0] input_423;
    input [0:0] input_424;
    input [0:0] input_425;
    input [0:0] input_426;
    input [0:0] input_427;
    input [0:0] input_428;
    input [0:0] input_429;
    input [0:0] input_430;
    input [0:0] input_431;
    input [0:0] input_432;
    input [0:0] input_433;
    input [0:0] input_434;
    input [0:0] input_435;
    input [0:0] input_436;
    input [0:0] input_437;
    input [0:0] input_438;
    input [0:0] input_439;
    input [0:0] input_440;
    input [0:0] input_441;
    input [0:0] input_442;
    input [0:0] input_443;
    input [0:0] input_444;
    input [0:0] input_445;
    input [0:0] input_446;
    input [0:0] input_447;
    input [0:0] input_448;
    input [0:0] input_449;
    input [0:0] input_450;
    input [0:0] input_451;
    input [0:0] input_452;
    input [0:0] input_453;
    input [0:0] input_454;
    input [0:0] input_455;
    input [0:0] input_456;
    input [0:0] input_457;
    input [0:0] input_458;
    input [0:0] input_459;
    input [0:0] input_460;
    input [0:0] input_461;
    input [0:0] input_462;
    input [0:0] input_463;
    input [0:0] input_464;
    input [0:0] input_465;
    input [0:0] input_466;
    input [0:0] input_467;
    input [0:0] input_468;
    input [0:0] input_469;
    input [0:0] input_470;
    input [0:0] input_471;
    input [0:0] input_472;
    input [0:0] input_473;
    input [0:0] input_474;
    input [0:0] input_475;
    input [0:0] input_476;
    input [0:0] input_477;
    input [0:0] input_478;
    input [0:0] input_479;
    input [0:0] input_480;
    input [0:0] input_481;
    input [0:0] input_482;
    input [0:0] input_483;
    input [0:0] input_484;
    input [0:0] input_485;
    input [0:0] input_486;
    input [0:0] input_487;
    input [0:0] input_488;
    input [0:0] input_489;
    input [0:0] input_490;
    input [0:0] input_491;
    input [0:0] input_492;
    input [0:0] input_493;
    input [0:0] input_494;
    input [0:0] input_495;
    input [0:0] input_496;
    input [0:0] input_497;
    input [0:0] input_498;
    input [0:0] input_499;
    input [0:0] input_500;
    input [0:0] input_501;
    input [0:0] input_502;
    input [0:0] input_503;
    input [0:0] input_504;
    input [0:0] input_505;
    input [0:0] input_506;
    input [0:0] input_507;
    input [0:0] input_508;
    input [0:0] input_509;
    input [0:0] input_510;
    input [0:0] input_511;
    input [0:0] input_512;
    input [0:0] input_513;
    input [0:0] input_514;
    input [0:0] input_515;
    input [0:0] input_516;
    input [0:0] input_517;
    input [0:0] input_518;
    input [0:0] input_519;
    input [0:0] input_520;
    input [0:0] input_521;
    input [0:0] input_522;
    input [0:0] input_523;
    input [0:0] input_524;
    input [0:0] input_525;
    input [0:0] input_526;
    input [0:0] input_527;
    input [0:0] input_528;
    input [0:0] input_529;
    input [0:0] input_530;
    input [0:0] input_531;
    input [0:0] input_532;
    input [0:0] input_533;
    input [0:0] input_534;
    input [0:0] input_535;
    input [0:0] input_536;
    input [0:0] input_537;
    input [0:0] input_538;
    input [0:0] input_539;
    input [0:0] input_540;
    input [0:0] input_541;
    input [0:0] input_542;
    input [0:0] input_543;
    input [0:0] input_544;
    input [0:0] input_545;
    input [0:0] input_546;
    input [0:0] input_547;
    input [0:0] input_548;
    input [0:0] input_549;
    input [0:0] input_550;
    input [0:0] input_551;
    input [0:0] input_552;
    input [0:0] input_553;
    input [0:0] input_554;
    input [0:0] input_555;
    input [0:0] input_556;
    input [0:0] input_557;
    input [0:0] input_558;
    input [0:0] input_559;
    input [0:0] input_560;
    input [0:0] input_561;
    input [0:0] input_562;
    input [0:0] input_563;
    input [0:0] input_564;
    input [0:0] input_565;
    input [0:0] input_566;
    input [0:0] input_567;
    input [0:0] input_568;
    input [0:0] input_569;
    input [0:0] input_570;
    input [0:0] input_571;
    input [0:0] input_572;
    input [0:0] input_573;
    input [0:0] input_574;
    input [0:0] input_575;
    input [0:0] input_576;
    input [0:0] input_577;
    input [0:0] input_578;
    input [0:0] input_579;
    input [0:0] input_580;
    input [0:0] input_581;
    input [0:0] input_582;
    input [0:0] input_583;
    input [0:0] input_584;
    input [0:0] input_585;
    input [0:0] input_586;
    input [0:0] input_587;
    input [0:0] input_588;
    input [0:0] input_589;
    input [0:0] input_590;
    input [0:0] input_591;
    input [0:0] input_592;
    input [0:0] input_593;
    input [0:0] input_594;
    input [0:0] input_595;
    input [0:0] input_596;
    input [0:0] input_597;
    input [0:0] input_598;
    input [0:0] input_599;
    input [0:0] input_600;
    input [0:0] input_601;
    input [0:0] input_602;
    input [0:0] input_603;
    input [0:0] input_604;
    input [0:0] input_605;
    input [0:0] input_606;
    input [0:0] input_607;
    input [0:0] input_608;
    input [0:0] input_609;
    input [0:0] input_610;
    input [0:0] input_611;
    input [0:0] input_612;
    input [0:0] input_613;
    input [0:0] input_614;
    input [0:0] input_615;
    input [0:0] input_616;
    input [0:0] input_617;
    input [0:0] input_618;
    input [0:0] input_619;
    input [0:0] input_620;
    input [0:0] input_621;
    input [0:0] input_622;
    input [0:0] input_623;
    input [0:0] input_624;
    input [0:0] input_625;
    input [0:0] input_626;
    input [0:0] input_627;
    input [0:0] input_628;
    input [0:0] input_629;
    input [0:0] input_630;
    input [0:0] input_631;
    input [0:0] input_632;
    input [0:0] input_633;
    input [0:0] input_634;
    input [0:0] input_635;
    input [0:0] input_636;
    input [0:0] input_637;
    input [0:0] input_638;
    input [0:0] input_639;
    input [0:0] input_640;
    input [0:0] input_641;
    input [0:0] input_642;
    input [0:0] input_643;
    input [0:0] input_644;
    input [0:0] input_645;
    input [0:0] input_646;
    input [0:0] input_647;
    input [0:0] input_648;
    input [0:0] input_649;
    input [0:0] input_650;
    input [0:0] input_651;
    input [0:0] input_652;
    input [0:0] input_653;
    input [0:0] input_654;
    input [0:0] input_655;
    input [0:0] input_656;
    input [0:0] input_657;
    input [0:0] input_658;
    input [0:0] input_659;
    input [0:0] input_660;
    input [0:0] input_661;
    input [0:0] input_662;
    input [0:0] input_663;
    input [0:0] input_664;
    input [0:0] input_665;
    input [0:0] input_666;
    input [0:0] input_667;
    input [0:0] input_668;
    input [0:0] input_669;
    input [0:0] input_670;
    input [0:0] input_671;
    input [0:0] input_672;
    input [0:0] input_673;
    input [0:0] input_674;
    input [0:0] input_675;
    input [0:0] input_676;
    input [0:0] input_677;
    input [0:0] input_678;
    input [0:0] input_679;
    input [0:0] input_680;
    input [0:0] input_681;
    input [0:0] input_682;
    input [0:0] input_683;
    input [0:0] input_684;
    input [0:0] input_685;
    input [0:0] input_686;
    input [0:0] input_687;
    input [0:0] input_688;
    input [0:0] input_689;
    input [0:0] input_690;
    input [0:0] input_691;
    input [0:0] input_692;
    input [0:0] input_693;
    input [0:0] input_694;
    input [0:0] input_695;
    input [0:0] input_696;
    input [0:0] input_697;
    input [0:0] input_698;
    input [0:0] input_699;
    input [0:0] input_700;
    input [0:0] input_701;
    input [0:0] input_702;
    input [0:0] input_703;
    input [0:0] input_704;
    input [0:0] input_705;
    input [0:0] input_706;
    input [0:0] input_707;
    input [0:0] input_708;
    input [0:0] input_709;
    input [0:0] input_710;
    input [0:0] input_711;
    input [0:0] input_712;
    input [0:0] input_713;
    input [0:0] input_714;
    input [0:0] input_715;
    input [0:0] input_716;
    input [0:0] input_717;
    input [0:0] input_718;
    input [0:0] input_719;
    input [0:0] input_720;
    input [0:0] input_721;
    input [0:0] input_722;
    input [0:0] input_723;
    input [0:0] input_724;
    input [0:0] input_725;
    input [0:0] input_726;
    input [0:0] input_727;
    input [0:0] input_728;
    input [0:0] input_729;
    input [0:0] input_730;
    input [0:0] input_731;
    input [0:0] input_732;
    input [0:0] input_733;
    input [0:0] input_734;
    input [0:0] input_735;
    input [0:0] input_736;
    input [0:0] input_737;
    input [0:0] input_738;
    input [0:0] input_739;
    input [0:0] input_740;
    input [0:0] input_741;
    input [0:0] input_742;
    input [0:0] input_743;
    input [0:0] input_744;
    input [0:0] input_745;
    input [0:0] input_746;
    input [0:0] input_747;
    input [0:0] input_748;
    input [0:0] input_749;
    input [0:0] input_750;
    input [0:0] input_751;
    input [0:0] input_752;
    input [0:0] input_753;
    input [0:0] input_754;
    input [0:0] input_755;
    input [0:0] input_756;
    input [0:0] input_757;
    input [0:0] input_758;
    input [0:0] input_759;
    input [0:0] input_760;
    input [0:0] input_761;
    input [0:0] input_762;
    input [0:0] input_763;
    input [0:0] input_764;
    input [0:0] input_765;
    input [0:0] input_766;
    input [0:0] input_767;
    input [0:0] input_768;
    input [0:0] input_769;
    input [0:0] input_770;
    input [0:0] input_771;
    input [0:0] input_772;
    input [0:0] input_773;
    input [0:0] input_774;
    input [0:0] input_775;
    input [0:0] input_776;
    input [0:0] input_777;
    input [0:0] input_778;
    input [0:0] input_779;
    input [0:0] input_780;
    input [0:0] input_781;
    input [0:0] input_782;
    input [0:0] input_783;
    input [0:0] input_784;
    input [0:0] input_785;
    input [0:0] input_786;
    input [0:0] input_787;
    input [0:0] input_788;
    input [0:0] input_789;
    input [0:0] input_790;
    input [0:0] input_791;
    input [0:0] input_792;
    input [0:0] input_793;
    input [0:0] input_794;
    input [0:0] input_795;
    input [0:0] input_796;
    input [0:0] input_797;
    input [0:0] input_798;
    input [0:0] input_799;
    input [0:0] input_800;
    input [0:0] input_801;
    input [0:0] input_802;
    input [0:0] input_803;
    input [0:0] input_804;
    input [0:0] input_805;
    input [0:0] input_806;
    input [0:0] input_807;
    input [0:0] input_808;
    input [0:0] input_809;
    input [0:0] input_810;
    input [0:0] input_811;
    input [0:0] input_812;
    input [0:0] input_813;
    input [0:0] input_814;
    input [0:0] input_815;
    input [0:0] input_816;
    input [0:0] input_817;
    input [0:0] input_818;
    input [0:0] input_819;
    input [0:0] input_820;
    input [0:0] input_821;
    input [0:0] input_822;
    input [0:0] input_823;
    input [0:0] input_824;
    input [0:0] input_825;
    input [0:0] input_826;
    input [0:0] input_827;
    input [0:0] input_828;
    input [0:0] input_829;
    input [0:0] input_830;
    input [0:0] input_831;
    input [0:0] input_832;
    input [0:0] input_833;
    input [0:0] input_834;
    input [0:0] input_835;
    input [0:0] input_836;
    input [0:0] input_837;
    input [0:0] input_838;
    input [0:0] input_839;
    input [0:0] input_840;
    input [0:0] input_841;
    input [0:0] input_842;
    input [0:0] input_843;
    input [0:0] input_844;
    input [0:0] input_845;
    input [0:0] input_846;
    input [0:0] input_847;
    input [0:0] input_848;
    input [0:0] input_849;
    input [0:0] input_850;
    input [0:0] input_851;
    input [0:0] input_852;
    input [0:0] input_853;
    input [0:0] input_854;
    input [0:0] input_855;
    input [0:0] input_856;
    input [0:0] input_857;
    input [0:0] input_858;
    input [0:0] input_859;
    input [0:0] input_860;
    input [0:0] input_861;
    input [0:0] input_862;
    input [0:0] input_863;
    input [0:0] input_864;
    input [0:0] input_865;
    input [0:0] input_866;
    input [0:0] input_867;
    input [0:0] input_868;
    input [0:0] input_869;
    input [0:0] input_870;
    input [0:0] input_871;
    input [0:0] input_872;
    input [0:0] input_873;
    input [0:0] input_874;
    input [0:0] input_875;
    input [0:0] input_876;
    input [0:0] input_877;
    input [0:0] input_878;
    input [0:0] input_879;
    input [0:0] input_880;
    input [0:0] input_881;
    input [0:0] input_882;
    input [0:0] input_883;
    input [0:0] input_884;
    input [0:0] input_885;
    input [0:0] input_886;
    input [0:0] input_887;
    input [0:0] input_888;
    input [0:0] input_889;
    input [0:0] input_890;
    input [0:0] input_891;
    input [0:0] input_892;
    input [0:0] input_893;
    input [0:0] input_894;
    input [0:0] input_895;
    input [0:0] input_896;
    input [0:0] input_897;
    input [0:0] input_898;
    input [0:0] input_899;
    input [0:0] input_900;
    input [0:0] input_901;
    input [0:0] input_902;
    input [0:0] input_903;
    input [0:0] input_904;
    input [0:0] input_905;
    input [0:0] input_906;
    input [0:0] input_907;
    input [0:0] input_908;
    input [0:0] input_909;
    input [0:0] input_910;
    input [0:0] input_911;
    input [0:0] input_912;
    input [0:0] input_913;
    input [0:0] input_914;
    input [0:0] input_915;
    input [0:0] input_916;
    input [0:0] input_917;
    input [0:0] input_918;
    input [0:0] input_919;
    input [0:0] input_920;
    input [0:0] input_921;
    input [0:0] input_922;
    input [0:0] input_923;
    input [0:0] input_924;
    input [0:0] input_925;
    input [0:0] input_926;
    input [0:0] input_927;
    input [0:0] input_928;
    input [0:0] input_929;
    input [0:0] input_930;
    input [0:0] input_931;
    input [0:0] input_932;
    input [0:0] input_933;
    input [0:0] input_934;
    input [0:0] input_935;
    input [0:0] input_936;
    input [0:0] input_937;
    input [0:0] input_938;
    input [0:0] input_939;
    input [0:0] input_940;
    input [0:0] input_941;
    input [0:0] input_942;
    input [0:0] input_943;
    input [0:0] input_944;
    input [0:0] input_945;
    input [0:0] input_946;
    input [0:0] input_947;
    input [0:0] input_948;
    input [0:0] input_949;
    input [0:0] input_950;
    input [0:0] input_951;
    input [0:0] input_952;
    input [0:0] input_953;
    input [0:0] input_954;
    input [0:0] input_955;
    input [0:0] input_956;
    input [0:0] input_957;
    input [0:0] input_958;
    input [0:0] input_959;
    input [0:0] input_960;
    input [0:0] input_961;
    input [0:0] input_962;
    input [0:0] input_963;
    input [0:0] input_964;
    input [0:0] input_965;
    input [0:0] input_966;
    input [0:0] input_967;
    input [0:0] input_968;
    input [0:0] input_969;
    input [0:0] input_970;
    input [0:0] input_971;
    input [0:0] input_972;
    input [0:0] input_973;
    input [0:0] input_974;
    input [0:0] input_975;
    input [0:0] input_976;
    input [0:0] input_977;
    input [0:0] input_978;
    input [0:0] input_979;
    input [0:0] input_980;
    input [0:0] input_981;
    input [0:0] input_982;
    input [0:0] input_983;
    input [0:0] input_984;
    input [0:0] input_985;
    input [0:0] input_986;
    input [0:0] input_987;
    input [0:0] input_988;
    input [0:0] input_989;
    input [0:0] input_990;
    input [0:0] input_991;
    input [0:0] input_992;
    input [0:0] input_993;
    input [0:0] input_994;
    input [0:0] input_995;
    input [0:0] input_996;
    input [0:0] input_997;
    input [0:0] input_998;
    input [0:0] input_999;
    input [0:0] input_1000;
    input [0:0] input_1001;
    input [0:0] input_1002;
    input [0:0] input_1003;
    input [0:0] input_1004;
    input [0:0] input_1005;
    input [0:0] input_1006;
    input [0:0] input_1007;
    input [0:0] input_1008;
    input [0:0] input_1009;
    input [0:0] input_1010;
    input [0:0] input_1011;
    input [0:0] input_1012;
    input [0:0] input_1013;
    input [0:0] input_1014;
    input [0:0] input_1015;
    input [0:0] input_1016;
    input [0:0] input_1017;
    input [0:0] input_1018;
    input [0:0] input_1019;
    input [0:0] input_1020;
    input [0:0] input_1021;
    input [0:0] input_1022;
    input [0:0] input_1023;
    input [9:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      10'b0000000000 : begin
        result = input_0;
      end
      10'b0000000001 : begin
        result = input_1;
      end
      10'b0000000010 : begin
        result = input_2;
      end
      10'b0000000011 : begin
        result = input_3;
      end
      10'b0000000100 : begin
        result = input_4;
      end
      10'b0000000101 : begin
        result = input_5;
      end
      10'b0000000110 : begin
        result = input_6;
      end
      10'b0000000111 : begin
        result = input_7;
      end
      10'b0000001000 : begin
        result = input_8;
      end
      10'b0000001001 : begin
        result = input_9;
      end
      10'b0000001010 : begin
        result = input_10;
      end
      10'b0000001011 : begin
        result = input_11;
      end
      10'b0000001100 : begin
        result = input_12;
      end
      10'b0000001101 : begin
        result = input_13;
      end
      10'b0000001110 : begin
        result = input_14;
      end
      10'b0000001111 : begin
        result = input_15;
      end
      10'b0000010000 : begin
        result = input_16;
      end
      10'b0000010001 : begin
        result = input_17;
      end
      10'b0000010010 : begin
        result = input_18;
      end
      10'b0000010011 : begin
        result = input_19;
      end
      10'b0000010100 : begin
        result = input_20;
      end
      10'b0000010101 : begin
        result = input_21;
      end
      10'b0000010110 : begin
        result = input_22;
      end
      10'b0000010111 : begin
        result = input_23;
      end
      10'b0000011000 : begin
        result = input_24;
      end
      10'b0000011001 : begin
        result = input_25;
      end
      10'b0000011010 : begin
        result = input_26;
      end
      10'b0000011011 : begin
        result = input_27;
      end
      10'b0000011100 : begin
        result = input_28;
      end
      10'b0000011101 : begin
        result = input_29;
      end
      10'b0000011110 : begin
        result = input_30;
      end
      10'b0000011111 : begin
        result = input_31;
      end
      10'b0000100000 : begin
        result = input_32;
      end
      10'b0000100001 : begin
        result = input_33;
      end
      10'b0000100010 : begin
        result = input_34;
      end
      10'b0000100011 : begin
        result = input_35;
      end
      10'b0000100100 : begin
        result = input_36;
      end
      10'b0000100101 : begin
        result = input_37;
      end
      10'b0000100110 : begin
        result = input_38;
      end
      10'b0000100111 : begin
        result = input_39;
      end
      10'b0000101000 : begin
        result = input_40;
      end
      10'b0000101001 : begin
        result = input_41;
      end
      10'b0000101010 : begin
        result = input_42;
      end
      10'b0000101011 : begin
        result = input_43;
      end
      10'b0000101100 : begin
        result = input_44;
      end
      10'b0000101101 : begin
        result = input_45;
      end
      10'b0000101110 : begin
        result = input_46;
      end
      10'b0000101111 : begin
        result = input_47;
      end
      10'b0000110000 : begin
        result = input_48;
      end
      10'b0000110001 : begin
        result = input_49;
      end
      10'b0000110010 : begin
        result = input_50;
      end
      10'b0000110011 : begin
        result = input_51;
      end
      10'b0000110100 : begin
        result = input_52;
      end
      10'b0000110101 : begin
        result = input_53;
      end
      10'b0000110110 : begin
        result = input_54;
      end
      10'b0000110111 : begin
        result = input_55;
      end
      10'b0000111000 : begin
        result = input_56;
      end
      10'b0000111001 : begin
        result = input_57;
      end
      10'b0000111010 : begin
        result = input_58;
      end
      10'b0000111011 : begin
        result = input_59;
      end
      10'b0000111100 : begin
        result = input_60;
      end
      10'b0000111101 : begin
        result = input_61;
      end
      10'b0000111110 : begin
        result = input_62;
      end
      10'b0000111111 : begin
        result = input_63;
      end
      10'b0001000000 : begin
        result = input_64;
      end
      10'b0001000001 : begin
        result = input_65;
      end
      10'b0001000010 : begin
        result = input_66;
      end
      10'b0001000011 : begin
        result = input_67;
      end
      10'b0001000100 : begin
        result = input_68;
      end
      10'b0001000101 : begin
        result = input_69;
      end
      10'b0001000110 : begin
        result = input_70;
      end
      10'b0001000111 : begin
        result = input_71;
      end
      10'b0001001000 : begin
        result = input_72;
      end
      10'b0001001001 : begin
        result = input_73;
      end
      10'b0001001010 : begin
        result = input_74;
      end
      10'b0001001011 : begin
        result = input_75;
      end
      10'b0001001100 : begin
        result = input_76;
      end
      10'b0001001101 : begin
        result = input_77;
      end
      10'b0001001110 : begin
        result = input_78;
      end
      10'b0001001111 : begin
        result = input_79;
      end
      10'b0001010000 : begin
        result = input_80;
      end
      10'b0001010001 : begin
        result = input_81;
      end
      10'b0001010010 : begin
        result = input_82;
      end
      10'b0001010011 : begin
        result = input_83;
      end
      10'b0001010100 : begin
        result = input_84;
      end
      10'b0001010101 : begin
        result = input_85;
      end
      10'b0001010110 : begin
        result = input_86;
      end
      10'b0001010111 : begin
        result = input_87;
      end
      10'b0001011000 : begin
        result = input_88;
      end
      10'b0001011001 : begin
        result = input_89;
      end
      10'b0001011010 : begin
        result = input_90;
      end
      10'b0001011011 : begin
        result = input_91;
      end
      10'b0001011100 : begin
        result = input_92;
      end
      10'b0001011101 : begin
        result = input_93;
      end
      10'b0001011110 : begin
        result = input_94;
      end
      10'b0001011111 : begin
        result = input_95;
      end
      10'b0001100000 : begin
        result = input_96;
      end
      10'b0001100001 : begin
        result = input_97;
      end
      10'b0001100010 : begin
        result = input_98;
      end
      10'b0001100011 : begin
        result = input_99;
      end
      10'b0001100100 : begin
        result = input_100;
      end
      10'b0001100101 : begin
        result = input_101;
      end
      10'b0001100110 : begin
        result = input_102;
      end
      10'b0001100111 : begin
        result = input_103;
      end
      10'b0001101000 : begin
        result = input_104;
      end
      10'b0001101001 : begin
        result = input_105;
      end
      10'b0001101010 : begin
        result = input_106;
      end
      10'b0001101011 : begin
        result = input_107;
      end
      10'b0001101100 : begin
        result = input_108;
      end
      10'b0001101101 : begin
        result = input_109;
      end
      10'b0001101110 : begin
        result = input_110;
      end
      10'b0001101111 : begin
        result = input_111;
      end
      10'b0001110000 : begin
        result = input_112;
      end
      10'b0001110001 : begin
        result = input_113;
      end
      10'b0001110010 : begin
        result = input_114;
      end
      10'b0001110011 : begin
        result = input_115;
      end
      10'b0001110100 : begin
        result = input_116;
      end
      10'b0001110101 : begin
        result = input_117;
      end
      10'b0001110110 : begin
        result = input_118;
      end
      10'b0001110111 : begin
        result = input_119;
      end
      10'b0001111000 : begin
        result = input_120;
      end
      10'b0001111001 : begin
        result = input_121;
      end
      10'b0001111010 : begin
        result = input_122;
      end
      10'b0001111011 : begin
        result = input_123;
      end
      10'b0001111100 : begin
        result = input_124;
      end
      10'b0001111101 : begin
        result = input_125;
      end
      10'b0001111110 : begin
        result = input_126;
      end
      10'b0001111111 : begin
        result = input_127;
      end
      10'b0010000000 : begin
        result = input_128;
      end
      10'b0010000001 : begin
        result = input_129;
      end
      10'b0010000010 : begin
        result = input_130;
      end
      10'b0010000011 : begin
        result = input_131;
      end
      10'b0010000100 : begin
        result = input_132;
      end
      10'b0010000101 : begin
        result = input_133;
      end
      10'b0010000110 : begin
        result = input_134;
      end
      10'b0010000111 : begin
        result = input_135;
      end
      10'b0010001000 : begin
        result = input_136;
      end
      10'b0010001001 : begin
        result = input_137;
      end
      10'b0010001010 : begin
        result = input_138;
      end
      10'b0010001011 : begin
        result = input_139;
      end
      10'b0010001100 : begin
        result = input_140;
      end
      10'b0010001101 : begin
        result = input_141;
      end
      10'b0010001110 : begin
        result = input_142;
      end
      10'b0010001111 : begin
        result = input_143;
      end
      10'b0010010000 : begin
        result = input_144;
      end
      10'b0010010001 : begin
        result = input_145;
      end
      10'b0010010010 : begin
        result = input_146;
      end
      10'b0010010011 : begin
        result = input_147;
      end
      10'b0010010100 : begin
        result = input_148;
      end
      10'b0010010101 : begin
        result = input_149;
      end
      10'b0010010110 : begin
        result = input_150;
      end
      10'b0010010111 : begin
        result = input_151;
      end
      10'b0010011000 : begin
        result = input_152;
      end
      10'b0010011001 : begin
        result = input_153;
      end
      10'b0010011010 : begin
        result = input_154;
      end
      10'b0010011011 : begin
        result = input_155;
      end
      10'b0010011100 : begin
        result = input_156;
      end
      10'b0010011101 : begin
        result = input_157;
      end
      10'b0010011110 : begin
        result = input_158;
      end
      10'b0010011111 : begin
        result = input_159;
      end
      10'b0010100000 : begin
        result = input_160;
      end
      10'b0010100001 : begin
        result = input_161;
      end
      10'b0010100010 : begin
        result = input_162;
      end
      10'b0010100011 : begin
        result = input_163;
      end
      10'b0010100100 : begin
        result = input_164;
      end
      10'b0010100101 : begin
        result = input_165;
      end
      10'b0010100110 : begin
        result = input_166;
      end
      10'b0010100111 : begin
        result = input_167;
      end
      10'b0010101000 : begin
        result = input_168;
      end
      10'b0010101001 : begin
        result = input_169;
      end
      10'b0010101010 : begin
        result = input_170;
      end
      10'b0010101011 : begin
        result = input_171;
      end
      10'b0010101100 : begin
        result = input_172;
      end
      10'b0010101101 : begin
        result = input_173;
      end
      10'b0010101110 : begin
        result = input_174;
      end
      10'b0010101111 : begin
        result = input_175;
      end
      10'b0010110000 : begin
        result = input_176;
      end
      10'b0010110001 : begin
        result = input_177;
      end
      10'b0010110010 : begin
        result = input_178;
      end
      10'b0010110011 : begin
        result = input_179;
      end
      10'b0010110100 : begin
        result = input_180;
      end
      10'b0010110101 : begin
        result = input_181;
      end
      10'b0010110110 : begin
        result = input_182;
      end
      10'b0010110111 : begin
        result = input_183;
      end
      10'b0010111000 : begin
        result = input_184;
      end
      10'b0010111001 : begin
        result = input_185;
      end
      10'b0010111010 : begin
        result = input_186;
      end
      10'b0010111011 : begin
        result = input_187;
      end
      10'b0010111100 : begin
        result = input_188;
      end
      10'b0010111101 : begin
        result = input_189;
      end
      10'b0010111110 : begin
        result = input_190;
      end
      10'b0010111111 : begin
        result = input_191;
      end
      10'b0011000000 : begin
        result = input_192;
      end
      10'b0011000001 : begin
        result = input_193;
      end
      10'b0011000010 : begin
        result = input_194;
      end
      10'b0011000011 : begin
        result = input_195;
      end
      10'b0011000100 : begin
        result = input_196;
      end
      10'b0011000101 : begin
        result = input_197;
      end
      10'b0011000110 : begin
        result = input_198;
      end
      10'b0011000111 : begin
        result = input_199;
      end
      10'b0011001000 : begin
        result = input_200;
      end
      10'b0011001001 : begin
        result = input_201;
      end
      10'b0011001010 : begin
        result = input_202;
      end
      10'b0011001011 : begin
        result = input_203;
      end
      10'b0011001100 : begin
        result = input_204;
      end
      10'b0011001101 : begin
        result = input_205;
      end
      10'b0011001110 : begin
        result = input_206;
      end
      10'b0011001111 : begin
        result = input_207;
      end
      10'b0011010000 : begin
        result = input_208;
      end
      10'b0011010001 : begin
        result = input_209;
      end
      10'b0011010010 : begin
        result = input_210;
      end
      10'b0011010011 : begin
        result = input_211;
      end
      10'b0011010100 : begin
        result = input_212;
      end
      10'b0011010101 : begin
        result = input_213;
      end
      10'b0011010110 : begin
        result = input_214;
      end
      10'b0011010111 : begin
        result = input_215;
      end
      10'b0011011000 : begin
        result = input_216;
      end
      10'b0011011001 : begin
        result = input_217;
      end
      10'b0011011010 : begin
        result = input_218;
      end
      10'b0011011011 : begin
        result = input_219;
      end
      10'b0011011100 : begin
        result = input_220;
      end
      10'b0011011101 : begin
        result = input_221;
      end
      10'b0011011110 : begin
        result = input_222;
      end
      10'b0011011111 : begin
        result = input_223;
      end
      10'b0011100000 : begin
        result = input_224;
      end
      10'b0011100001 : begin
        result = input_225;
      end
      10'b0011100010 : begin
        result = input_226;
      end
      10'b0011100011 : begin
        result = input_227;
      end
      10'b0011100100 : begin
        result = input_228;
      end
      10'b0011100101 : begin
        result = input_229;
      end
      10'b0011100110 : begin
        result = input_230;
      end
      10'b0011100111 : begin
        result = input_231;
      end
      10'b0011101000 : begin
        result = input_232;
      end
      10'b0011101001 : begin
        result = input_233;
      end
      10'b0011101010 : begin
        result = input_234;
      end
      10'b0011101011 : begin
        result = input_235;
      end
      10'b0011101100 : begin
        result = input_236;
      end
      10'b0011101101 : begin
        result = input_237;
      end
      10'b0011101110 : begin
        result = input_238;
      end
      10'b0011101111 : begin
        result = input_239;
      end
      10'b0011110000 : begin
        result = input_240;
      end
      10'b0011110001 : begin
        result = input_241;
      end
      10'b0011110010 : begin
        result = input_242;
      end
      10'b0011110011 : begin
        result = input_243;
      end
      10'b0011110100 : begin
        result = input_244;
      end
      10'b0011110101 : begin
        result = input_245;
      end
      10'b0011110110 : begin
        result = input_246;
      end
      10'b0011110111 : begin
        result = input_247;
      end
      10'b0011111000 : begin
        result = input_248;
      end
      10'b0011111001 : begin
        result = input_249;
      end
      10'b0011111010 : begin
        result = input_250;
      end
      10'b0011111011 : begin
        result = input_251;
      end
      10'b0011111100 : begin
        result = input_252;
      end
      10'b0011111101 : begin
        result = input_253;
      end
      10'b0011111110 : begin
        result = input_254;
      end
      10'b0011111111 : begin
        result = input_255;
      end
      10'b0100000000 : begin
        result = input_256;
      end
      10'b0100000001 : begin
        result = input_257;
      end
      10'b0100000010 : begin
        result = input_258;
      end
      10'b0100000011 : begin
        result = input_259;
      end
      10'b0100000100 : begin
        result = input_260;
      end
      10'b0100000101 : begin
        result = input_261;
      end
      10'b0100000110 : begin
        result = input_262;
      end
      10'b0100000111 : begin
        result = input_263;
      end
      10'b0100001000 : begin
        result = input_264;
      end
      10'b0100001001 : begin
        result = input_265;
      end
      10'b0100001010 : begin
        result = input_266;
      end
      10'b0100001011 : begin
        result = input_267;
      end
      10'b0100001100 : begin
        result = input_268;
      end
      10'b0100001101 : begin
        result = input_269;
      end
      10'b0100001110 : begin
        result = input_270;
      end
      10'b0100001111 : begin
        result = input_271;
      end
      10'b0100010000 : begin
        result = input_272;
      end
      10'b0100010001 : begin
        result = input_273;
      end
      10'b0100010010 : begin
        result = input_274;
      end
      10'b0100010011 : begin
        result = input_275;
      end
      10'b0100010100 : begin
        result = input_276;
      end
      10'b0100010101 : begin
        result = input_277;
      end
      10'b0100010110 : begin
        result = input_278;
      end
      10'b0100010111 : begin
        result = input_279;
      end
      10'b0100011000 : begin
        result = input_280;
      end
      10'b0100011001 : begin
        result = input_281;
      end
      10'b0100011010 : begin
        result = input_282;
      end
      10'b0100011011 : begin
        result = input_283;
      end
      10'b0100011100 : begin
        result = input_284;
      end
      10'b0100011101 : begin
        result = input_285;
      end
      10'b0100011110 : begin
        result = input_286;
      end
      10'b0100011111 : begin
        result = input_287;
      end
      10'b0100100000 : begin
        result = input_288;
      end
      10'b0100100001 : begin
        result = input_289;
      end
      10'b0100100010 : begin
        result = input_290;
      end
      10'b0100100011 : begin
        result = input_291;
      end
      10'b0100100100 : begin
        result = input_292;
      end
      10'b0100100101 : begin
        result = input_293;
      end
      10'b0100100110 : begin
        result = input_294;
      end
      10'b0100100111 : begin
        result = input_295;
      end
      10'b0100101000 : begin
        result = input_296;
      end
      10'b0100101001 : begin
        result = input_297;
      end
      10'b0100101010 : begin
        result = input_298;
      end
      10'b0100101011 : begin
        result = input_299;
      end
      10'b0100101100 : begin
        result = input_300;
      end
      10'b0100101101 : begin
        result = input_301;
      end
      10'b0100101110 : begin
        result = input_302;
      end
      10'b0100101111 : begin
        result = input_303;
      end
      10'b0100110000 : begin
        result = input_304;
      end
      10'b0100110001 : begin
        result = input_305;
      end
      10'b0100110010 : begin
        result = input_306;
      end
      10'b0100110011 : begin
        result = input_307;
      end
      10'b0100110100 : begin
        result = input_308;
      end
      10'b0100110101 : begin
        result = input_309;
      end
      10'b0100110110 : begin
        result = input_310;
      end
      10'b0100110111 : begin
        result = input_311;
      end
      10'b0100111000 : begin
        result = input_312;
      end
      10'b0100111001 : begin
        result = input_313;
      end
      10'b0100111010 : begin
        result = input_314;
      end
      10'b0100111011 : begin
        result = input_315;
      end
      10'b0100111100 : begin
        result = input_316;
      end
      10'b0100111101 : begin
        result = input_317;
      end
      10'b0100111110 : begin
        result = input_318;
      end
      10'b0100111111 : begin
        result = input_319;
      end
      10'b0101000000 : begin
        result = input_320;
      end
      10'b0101000001 : begin
        result = input_321;
      end
      10'b0101000010 : begin
        result = input_322;
      end
      10'b0101000011 : begin
        result = input_323;
      end
      10'b0101000100 : begin
        result = input_324;
      end
      10'b0101000101 : begin
        result = input_325;
      end
      10'b0101000110 : begin
        result = input_326;
      end
      10'b0101000111 : begin
        result = input_327;
      end
      10'b0101001000 : begin
        result = input_328;
      end
      10'b0101001001 : begin
        result = input_329;
      end
      10'b0101001010 : begin
        result = input_330;
      end
      10'b0101001011 : begin
        result = input_331;
      end
      10'b0101001100 : begin
        result = input_332;
      end
      10'b0101001101 : begin
        result = input_333;
      end
      10'b0101001110 : begin
        result = input_334;
      end
      10'b0101001111 : begin
        result = input_335;
      end
      10'b0101010000 : begin
        result = input_336;
      end
      10'b0101010001 : begin
        result = input_337;
      end
      10'b0101010010 : begin
        result = input_338;
      end
      10'b0101010011 : begin
        result = input_339;
      end
      10'b0101010100 : begin
        result = input_340;
      end
      10'b0101010101 : begin
        result = input_341;
      end
      10'b0101010110 : begin
        result = input_342;
      end
      10'b0101010111 : begin
        result = input_343;
      end
      10'b0101011000 : begin
        result = input_344;
      end
      10'b0101011001 : begin
        result = input_345;
      end
      10'b0101011010 : begin
        result = input_346;
      end
      10'b0101011011 : begin
        result = input_347;
      end
      10'b0101011100 : begin
        result = input_348;
      end
      10'b0101011101 : begin
        result = input_349;
      end
      10'b0101011110 : begin
        result = input_350;
      end
      10'b0101011111 : begin
        result = input_351;
      end
      10'b0101100000 : begin
        result = input_352;
      end
      10'b0101100001 : begin
        result = input_353;
      end
      10'b0101100010 : begin
        result = input_354;
      end
      10'b0101100011 : begin
        result = input_355;
      end
      10'b0101100100 : begin
        result = input_356;
      end
      10'b0101100101 : begin
        result = input_357;
      end
      10'b0101100110 : begin
        result = input_358;
      end
      10'b0101100111 : begin
        result = input_359;
      end
      10'b0101101000 : begin
        result = input_360;
      end
      10'b0101101001 : begin
        result = input_361;
      end
      10'b0101101010 : begin
        result = input_362;
      end
      10'b0101101011 : begin
        result = input_363;
      end
      10'b0101101100 : begin
        result = input_364;
      end
      10'b0101101101 : begin
        result = input_365;
      end
      10'b0101101110 : begin
        result = input_366;
      end
      10'b0101101111 : begin
        result = input_367;
      end
      10'b0101110000 : begin
        result = input_368;
      end
      10'b0101110001 : begin
        result = input_369;
      end
      10'b0101110010 : begin
        result = input_370;
      end
      10'b0101110011 : begin
        result = input_371;
      end
      10'b0101110100 : begin
        result = input_372;
      end
      10'b0101110101 : begin
        result = input_373;
      end
      10'b0101110110 : begin
        result = input_374;
      end
      10'b0101110111 : begin
        result = input_375;
      end
      10'b0101111000 : begin
        result = input_376;
      end
      10'b0101111001 : begin
        result = input_377;
      end
      10'b0101111010 : begin
        result = input_378;
      end
      10'b0101111011 : begin
        result = input_379;
      end
      10'b0101111100 : begin
        result = input_380;
      end
      10'b0101111101 : begin
        result = input_381;
      end
      10'b0101111110 : begin
        result = input_382;
      end
      10'b0101111111 : begin
        result = input_383;
      end
      10'b0110000000 : begin
        result = input_384;
      end
      10'b0110000001 : begin
        result = input_385;
      end
      10'b0110000010 : begin
        result = input_386;
      end
      10'b0110000011 : begin
        result = input_387;
      end
      10'b0110000100 : begin
        result = input_388;
      end
      10'b0110000101 : begin
        result = input_389;
      end
      10'b0110000110 : begin
        result = input_390;
      end
      10'b0110000111 : begin
        result = input_391;
      end
      10'b0110001000 : begin
        result = input_392;
      end
      10'b0110001001 : begin
        result = input_393;
      end
      10'b0110001010 : begin
        result = input_394;
      end
      10'b0110001011 : begin
        result = input_395;
      end
      10'b0110001100 : begin
        result = input_396;
      end
      10'b0110001101 : begin
        result = input_397;
      end
      10'b0110001110 : begin
        result = input_398;
      end
      10'b0110001111 : begin
        result = input_399;
      end
      10'b0110010000 : begin
        result = input_400;
      end
      10'b0110010001 : begin
        result = input_401;
      end
      10'b0110010010 : begin
        result = input_402;
      end
      10'b0110010011 : begin
        result = input_403;
      end
      10'b0110010100 : begin
        result = input_404;
      end
      10'b0110010101 : begin
        result = input_405;
      end
      10'b0110010110 : begin
        result = input_406;
      end
      10'b0110010111 : begin
        result = input_407;
      end
      10'b0110011000 : begin
        result = input_408;
      end
      10'b0110011001 : begin
        result = input_409;
      end
      10'b0110011010 : begin
        result = input_410;
      end
      10'b0110011011 : begin
        result = input_411;
      end
      10'b0110011100 : begin
        result = input_412;
      end
      10'b0110011101 : begin
        result = input_413;
      end
      10'b0110011110 : begin
        result = input_414;
      end
      10'b0110011111 : begin
        result = input_415;
      end
      10'b0110100000 : begin
        result = input_416;
      end
      10'b0110100001 : begin
        result = input_417;
      end
      10'b0110100010 : begin
        result = input_418;
      end
      10'b0110100011 : begin
        result = input_419;
      end
      10'b0110100100 : begin
        result = input_420;
      end
      10'b0110100101 : begin
        result = input_421;
      end
      10'b0110100110 : begin
        result = input_422;
      end
      10'b0110100111 : begin
        result = input_423;
      end
      10'b0110101000 : begin
        result = input_424;
      end
      10'b0110101001 : begin
        result = input_425;
      end
      10'b0110101010 : begin
        result = input_426;
      end
      10'b0110101011 : begin
        result = input_427;
      end
      10'b0110101100 : begin
        result = input_428;
      end
      10'b0110101101 : begin
        result = input_429;
      end
      10'b0110101110 : begin
        result = input_430;
      end
      10'b0110101111 : begin
        result = input_431;
      end
      10'b0110110000 : begin
        result = input_432;
      end
      10'b0110110001 : begin
        result = input_433;
      end
      10'b0110110010 : begin
        result = input_434;
      end
      10'b0110110011 : begin
        result = input_435;
      end
      10'b0110110100 : begin
        result = input_436;
      end
      10'b0110110101 : begin
        result = input_437;
      end
      10'b0110110110 : begin
        result = input_438;
      end
      10'b0110110111 : begin
        result = input_439;
      end
      10'b0110111000 : begin
        result = input_440;
      end
      10'b0110111001 : begin
        result = input_441;
      end
      10'b0110111010 : begin
        result = input_442;
      end
      10'b0110111011 : begin
        result = input_443;
      end
      10'b0110111100 : begin
        result = input_444;
      end
      10'b0110111101 : begin
        result = input_445;
      end
      10'b0110111110 : begin
        result = input_446;
      end
      10'b0110111111 : begin
        result = input_447;
      end
      10'b0111000000 : begin
        result = input_448;
      end
      10'b0111000001 : begin
        result = input_449;
      end
      10'b0111000010 : begin
        result = input_450;
      end
      10'b0111000011 : begin
        result = input_451;
      end
      10'b0111000100 : begin
        result = input_452;
      end
      10'b0111000101 : begin
        result = input_453;
      end
      10'b0111000110 : begin
        result = input_454;
      end
      10'b0111000111 : begin
        result = input_455;
      end
      10'b0111001000 : begin
        result = input_456;
      end
      10'b0111001001 : begin
        result = input_457;
      end
      10'b0111001010 : begin
        result = input_458;
      end
      10'b0111001011 : begin
        result = input_459;
      end
      10'b0111001100 : begin
        result = input_460;
      end
      10'b0111001101 : begin
        result = input_461;
      end
      10'b0111001110 : begin
        result = input_462;
      end
      10'b0111001111 : begin
        result = input_463;
      end
      10'b0111010000 : begin
        result = input_464;
      end
      10'b0111010001 : begin
        result = input_465;
      end
      10'b0111010010 : begin
        result = input_466;
      end
      10'b0111010011 : begin
        result = input_467;
      end
      10'b0111010100 : begin
        result = input_468;
      end
      10'b0111010101 : begin
        result = input_469;
      end
      10'b0111010110 : begin
        result = input_470;
      end
      10'b0111010111 : begin
        result = input_471;
      end
      10'b0111011000 : begin
        result = input_472;
      end
      10'b0111011001 : begin
        result = input_473;
      end
      10'b0111011010 : begin
        result = input_474;
      end
      10'b0111011011 : begin
        result = input_475;
      end
      10'b0111011100 : begin
        result = input_476;
      end
      10'b0111011101 : begin
        result = input_477;
      end
      10'b0111011110 : begin
        result = input_478;
      end
      10'b0111011111 : begin
        result = input_479;
      end
      10'b0111100000 : begin
        result = input_480;
      end
      10'b0111100001 : begin
        result = input_481;
      end
      10'b0111100010 : begin
        result = input_482;
      end
      10'b0111100011 : begin
        result = input_483;
      end
      10'b0111100100 : begin
        result = input_484;
      end
      10'b0111100101 : begin
        result = input_485;
      end
      10'b0111100110 : begin
        result = input_486;
      end
      10'b0111100111 : begin
        result = input_487;
      end
      10'b0111101000 : begin
        result = input_488;
      end
      10'b0111101001 : begin
        result = input_489;
      end
      10'b0111101010 : begin
        result = input_490;
      end
      10'b0111101011 : begin
        result = input_491;
      end
      10'b0111101100 : begin
        result = input_492;
      end
      10'b0111101101 : begin
        result = input_493;
      end
      10'b0111101110 : begin
        result = input_494;
      end
      10'b0111101111 : begin
        result = input_495;
      end
      10'b0111110000 : begin
        result = input_496;
      end
      10'b0111110001 : begin
        result = input_497;
      end
      10'b0111110010 : begin
        result = input_498;
      end
      10'b0111110011 : begin
        result = input_499;
      end
      10'b0111110100 : begin
        result = input_500;
      end
      10'b0111110101 : begin
        result = input_501;
      end
      10'b0111110110 : begin
        result = input_502;
      end
      10'b0111110111 : begin
        result = input_503;
      end
      10'b0111111000 : begin
        result = input_504;
      end
      10'b0111111001 : begin
        result = input_505;
      end
      10'b0111111010 : begin
        result = input_506;
      end
      10'b0111111011 : begin
        result = input_507;
      end
      10'b0111111100 : begin
        result = input_508;
      end
      10'b0111111101 : begin
        result = input_509;
      end
      10'b0111111110 : begin
        result = input_510;
      end
      10'b0111111111 : begin
        result = input_511;
      end
      10'b1000000000 : begin
        result = input_512;
      end
      10'b1000000001 : begin
        result = input_513;
      end
      10'b1000000010 : begin
        result = input_514;
      end
      10'b1000000011 : begin
        result = input_515;
      end
      10'b1000000100 : begin
        result = input_516;
      end
      10'b1000000101 : begin
        result = input_517;
      end
      10'b1000000110 : begin
        result = input_518;
      end
      10'b1000000111 : begin
        result = input_519;
      end
      10'b1000001000 : begin
        result = input_520;
      end
      10'b1000001001 : begin
        result = input_521;
      end
      10'b1000001010 : begin
        result = input_522;
      end
      10'b1000001011 : begin
        result = input_523;
      end
      10'b1000001100 : begin
        result = input_524;
      end
      10'b1000001101 : begin
        result = input_525;
      end
      10'b1000001110 : begin
        result = input_526;
      end
      10'b1000001111 : begin
        result = input_527;
      end
      10'b1000010000 : begin
        result = input_528;
      end
      10'b1000010001 : begin
        result = input_529;
      end
      10'b1000010010 : begin
        result = input_530;
      end
      10'b1000010011 : begin
        result = input_531;
      end
      10'b1000010100 : begin
        result = input_532;
      end
      10'b1000010101 : begin
        result = input_533;
      end
      10'b1000010110 : begin
        result = input_534;
      end
      10'b1000010111 : begin
        result = input_535;
      end
      10'b1000011000 : begin
        result = input_536;
      end
      10'b1000011001 : begin
        result = input_537;
      end
      10'b1000011010 : begin
        result = input_538;
      end
      10'b1000011011 : begin
        result = input_539;
      end
      10'b1000011100 : begin
        result = input_540;
      end
      10'b1000011101 : begin
        result = input_541;
      end
      10'b1000011110 : begin
        result = input_542;
      end
      10'b1000011111 : begin
        result = input_543;
      end
      10'b1000100000 : begin
        result = input_544;
      end
      10'b1000100001 : begin
        result = input_545;
      end
      10'b1000100010 : begin
        result = input_546;
      end
      10'b1000100011 : begin
        result = input_547;
      end
      10'b1000100100 : begin
        result = input_548;
      end
      10'b1000100101 : begin
        result = input_549;
      end
      10'b1000100110 : begin
        result = input_550;
      end
      10'b1000100111 : begin
        result = input_551;
      end
      10'b1000101000 : begin
        result = input_552;
      end
      10'b1000101001 : begin
        result = input_553;
      end
      10'b1000101010 : begin
        result = input_554;
      end
      10'b1000101011 : begin
        result = input_555;
      end
      10'b1000101100 : begin
        result = input_556;
      end
      10'b1000101101 : begin
        result = input_557;
      end
      10'b1000101110 : begin
        result = input_558;
      end
      10'b1000101111 : begin
        result = input_559;
      end
      10'b1000110000 : begin
        result = input_560;
      end
      10'b1000110001 : begin
        result = input_561;
      end
      10'b1000110010 : begin
        result = input_562;
      end
      10'b1000110011 : begin
        result = input_563;
      end
      10'b1000110100 : begin
        result = input_564;
      end
      10'b1000110101 : begin
        result = input_565;
      end
      10'b1000110110 : begin
        result = input_566;
      end
      10'b1000110111 : begin
        result = input_567;
      end
      10'b1000111000 : begin
        result = input_568;
      end
      10'b1000111001 : begin
        result = input_569;
      end
      10'b1000111010 : begin
        result = input_570;
      end
      10'b1000111011 : begin
        result = input_571;
      end
      10'b1000111100 : begin
        result = input_572;
      end
      10'b1000111101 : begin
        result = input_573;
      end
      10'b1000111110 : begin
        result = input_574;
      end
      10'b1000111111 : begin
        result = input_575;
      end
      10'b1001000000 : begin
        result = input_576;
      end
      10'b1001000001 : begin
        result = input_577;
      end
      10'b1001000010 : begin
        result = input_578;
      end
      10'b1001000011 : begin
        result = input_579;
      end
      10'b1001000100 : begin
        result = input_580;
      end
      10'b1001000101 : begin
        result = input_581;
      end
      10'b1001000110 : begin
        result = input_582;
      end
      10'b1001000111 : begin
        result = input_583;
      end
      10'b1001001000 : begin
        result = input_584;
      end
      10'b1001001001 : begin
        result = input_585;
      end
      10'b1001001010 : begin
        result = input_586;
      end
      10'b1001001011 : begin
        result = input_587;
      end
      10'b1001001100 : begin
        result = input_588;
      end
      10'b1001001101 : begin
        result = input_589;
      end
      10'b1001001110 : begin
        result = input_590;
      end
      10'b1001001111 : begin
        result = input_591;
      end
      10'b1001010000 : begin
        result = input_592;
      end
      10'b1001010001 : begin
        result = input_593;
      end
      10'b1001010010 : begin
        result = input_594;
      end
      10'b1001010011 : begin
        result = input_595;
      end
      10'b1001010100 : begin
        result = input_596;
      end
      10'b1001010101 : begin
        result = input_597;
      end
      10'b1001010110 : begin
        result = input_598;
      end
      10'b1001010111 : begin
        result = input_599;
      end
      10'b1001011000 : begin
        result = input_600;
      end
      10'b1001011001 : begin
        result = input_601;
      end
      10'b1001011010 : begin
        result = input_602;
      end
      10'b1001011011 : begin
        result = input_603;
      end
      10'b1001011100 : begin
        result = input_604;
      end
      10'b1001011101 : begin
        result = input_605;
      end
      10'b1001011110 : begin
        result = input_606;
      end
      10'b1001011111 : begin
        result = input_607;
      end
      10'b1001100000 : begin
        result = input_608;
      end
      10'b1001100001 : begin
        result = input_609;
      end
      10'b1001100010 : begin
        result = input_610;
      end
      10'b1001100011 : begin
        result = input_611;
      end
      10'b1001100100 : begin
        result = input_612;
      end
      10'b1001100101 : begin
        result = input_613;
      end
      10'b1001100110 : begin
        result = input_614;
      end
      10'b1001100111 : begin
        result = input_615;
      end
      10'b1001101000 : begin
        result = input_616;
      end
      10'b1001101001 : begin
        result = input_617;
      end
      10'b1001101010 : begin
        result = input_618;
      end
      10'b1001101011 : begin
        result = input_619;
      end
      10'b1001101100 : begin
        result = input_620;
      end
      10'b1001101101 : begin
        result = input_621;
      end
      10'b1001101110 : begin
        result = input_622;
      end
      10'b1001101111 : begin
        result = input_623;
      end
      10'b1001110000 : begin
        result = input_624;
      end
      10'b1001110001 : begin
        result = input_625;
      end
      10'b1001110010 : begin
        result = input_626;
      end
      10'b1001110011 : begin
        result = input_627;
      end
      10'b1001110100 : begin
        result = input_628;
      end
      10'b1001110101 : begin
        result = input_629;
      end
      10'b1001110110 : begin
        result = input_630;
      end
      10'b1001110111 : begin
        result = input_631;
      end
      10'b1001111000 : begin
        result = input_632;
      end
      10'b1001111001 : begin
        result = input_633;
      end
      10'b1001111010 : begin
        result = input_634;
      end
      10'b1001111011 : begin
        result = input_635;
      end
      10'b1001111100 : begin
        result = input_636;
      end
      10'b1001111101 : begin
        result = input_637;
      end
      10'b1001111110 : begin
        result = input_638;
      end
      10'b1001111111 : begin
        result = input_639;
      end
      10'b1010000000 : begin
        result = input_640;
      end
      10'b1010000001 : begin
        result = input_641;
      end
      10'b1010000010 : begin
        result = input_642;
      end
      10'b1010000011 : begin
        result = input_643;
      end
      10'b1010000100 : begin
        result = input_644;
      end
      10'b1010000101 : begin
        result = input_645;
      end
      10'b1010000110 : begin
        result = input_646;
      end
      10'b1010000111 : begin
        result = input_647;
      end
      10'b1010001000 : begin
        result = input_648;
      end
      10'b1010001001 : begin
        result = input_649;
      end
      10'b1010001010 : begin
        result = input_650;
      end
      10'b1010001011 : begin
        result = input_651;
      end
      10'b1010001100 : begin
        result = input_652;
      end
      10'b1010001101 : begin
        result = input_653;
      end
      10'b1010001110 : begin
        result = input_654;
      end
      10'b1010001111 : begin
        result = input_655;
      end
      10'b1010010000 : begin
        result = input_656;
      end
      10'b1010010001 : begin
        result = input_657;
      end
      10'b1010010010 : begin
        result = input_658;
      end
      10'b1010010011 : begin
        result = input_659;
      end
      10'b1010010100 : begin
        result = input_660;
      end
      10'b1010010101 : begin
        result = input_661;
      end
      10'b1010010110 : begin
        result = input_662;
      end
      10'b1010010111 : begin
        result = input_663;
      end
      10'b1010011000 : begin
        result = input_664;
      end
      10'b1010011001 : begin
        result = input_665;
      end
      10'b1010011010 : begin
        result = input_666;
      end
      10'b1010011011 : begin
        result = input_667;
      end
      10'b1010011100 : begin
        result = input_668;
      end
      10'b1010011101 : begin
        result = input_669;
      end
      10'b1010011110 : begin
        result = input_670;
      end
      10'b1010011111 : begin
        result = input_671;
      end
      10'b1010100000 : begin
        result = input_672;
      end
      10'b1010100001 : begin
        result = input_673;
      end
      10'b1010100010 : begin
        result = input_674;
      end
      10'b1010100011 : begin
        result = input_675;
      end
      10'b1010100100 : begin
        result = input_676;
      end
      10'b1010100101 : begin
        result = input_677;
      end
      10'b1010100110 : begin
        result = input_678;
      end
      10'b1010100111 : begin
        result = input_679;
      end
      10'b1010101000 : begin
        result = input_680;
      end
      10'b1010101001 : begin
        result = input_681;
      end
      10'b1010101010 : begin
        result = input_682;
      end
      10'b1010101011 : begin
        result = input_683;
      end
      10'b1010101100 : begin
        result = input_684;
      end
      10'b1010101101 : begin
        result = input_685;
      end
      10'b1010101110 : begin
        result = input_686;
      end
      10'b1010101111 : begin
        result = input_687;
      end
      10'b1010110000 : begin
        result = input_688;
      end
      10'b1010110001 : begin
        result = input_689;
      end
      10'b1010110010 : begin
        result = input_690;
      end
      10'b1010110011 : begin
        result = input_691;
      end
      10'b1010110100 : begin
        result = input_692;
      end
      10'b1010110101 : begin
        result = input_693;
      end
      10'b1010110110 : begin
        result = input_694;
      end
      10'b1010110111 : begin
        result = input_695;
      end
      10'b1010111000 : begin
        result = input_696;
      end
      10'b1010111001 : begin
        result = input_697;
      end
      10'b1010111010 : begin
        result = input_698;
      end
      10'b1010111011 : begin
        result = input_699;
      end
      10'b1010111100 : begin
        result = input_700;
      end
      10'b1010111101 : begin
        result = input_701;
      end
      10'b1010111110 : begin
        result = input_702;
      end
      10'b1010111111 : begin
        result = input_703;
      end
      10'b1011000000 : begin
        result = input_704;
      end
      10'b1011000001 : begin
        result = input_705;
      end
      10'b1011000010 : begin
        result = input_706;
      end
      10'b1011000011 : begin
        result = input_707;
      end
      10'b1011000100 : begin
        result = input_708;
      end
      10'b1011000101 : begin
        result = input_709;
      end
      10'b1011000110 : begin
        result = input_710;
      end
      10'b1011000111 : begin
        result = input_711;
      end
      10'b1011001000 : begin
        result = input_712;
      end
      10'b1011001001 : begin
        result = input_713;
      end
      10'b1011001010 : begin
        result = input_714;
      end
      10'b1011001011 : begin
        result = input_715;
      end
      10'b1011001100 : begin
        result = input_716;
      end
      10'b1011001101 : begin
        result = input_717;
      end
      10'b1011001110 : begin
        result = input_718;
      end
      10'b1011001111 : begin
        result = input_719;
      end
      10'b1011010000 : begin
        result = input_720;
      end
      10'b1011010001 : begin
        result = input_721;
      end
      10'b1011010010 : begin
        result = input_722;
      end
      10'b1011010011 : begin
        result = input_723;
      end
      10'b1011010100 : begin
        result = input_724;
      end
      10'b1011010101 : begin
        result = input_725;
      end
      10'b1011010110 : begin
        result = input_726;
      end
      10'b1011010111 : begin
        result = input_727;
      end
      10'b1011011000 : begin
        result = input_728;
      end
      10'b1011011001 : begin
        result = input_729;
      end
      10'b1011011010 : begin
        result = input_730;
      end
      10'b1011011011 : begin
        result = input_731;
      end
      10'b1011011100 : begin
        result = input_732;
      end
      10'b1011011101 : begin
        result = input_733;
      end
      10'b1011011110 : begin
        result = input_734;
      end
      10'b1011011111 : begin
        result = input_735;
      end
      10'b1011100000 : begin
        result = input_736;
      end
      10'b1011100001 : begin
        result = input_737;
      end
      10'b1011100010 : begin
        result = input_738;
      end
      10'b1011100011 : begin
        result = input_739;
      end
      10'b1011100100 : begin
        result = input_740;
      end
      10'b1011100101 : begin
        result = input_741;
      end
      10'b1011100110 : begin
        result = input_742;
      end
      10'b1011100111 : begin
        result = input_743;
      end
      10'b1011101000 : begin
        result = input_744;
      end
      10'b1011101001 : begin
        result = input_745;
      end
      10'b1011101010 : begin
        result = input_746;
      end
      10'b1011101011 : begin
        result = input_747;
      end
      10'b1011101100 : begin
        result = input_748;
      end
      10'b1011101101 : begin
        result = input_749;
      end
      10'b1011101110 : begin
        result = input_750;
      end
      10'b1011101111 : begin
        result = input_751;
      end
      10'b1011110000 : begin
        result = input_752;
      end
      10'b1011110001 : begin
        result = input_753;
      end
      10'b1011110010 : begin
        result = input_754;
      end
      10'b1011110011 : begin
        result = input_755;
      end
      10'b1011110100 : begin
        result = input_756;
      end
      10'b1011110101 : begin
        result = input_757;
      end
      10'b1011110110 : begin
        result = input_758;
      end
      10'b1011110111 : begin
        result = input_759;
      end
      10'b1011111000 : begin
        result = input_760;
      end
      10'b1011111001 : begin
        result = input_761;
      end
      10'b1011111010 : begin
        result = input_762;
      end
      10'b1011111011 : begin
        result = input_763;
      end
      10'b1011111100 : begin
        result = input_764;
      end
      10'b1011111101 : begin
        result = input_765;
      end
      10'b1011111110 : begin
        result = input_766;
      end
      10'b1011111111 : begin
        result = input_767;
      end
      10'b1100000000 : begin
        result = input_768;
      end
      10'b1100000001 : begin
        result = input_769;
      end
      10'b1100000010 : begin
        result = input_770;
      end
      10'b1100000011 : begin
        result = input_771;
      end
      10'b1100000100 : begin
        result = input_772;
      end
      10'b1100000101 : begin
        result = input_773;
      end
      10'b1100000110 : begin
        result = input_774;
      end
      10'b1100000111 : begin
        result = input_775;
      end
      10'b1100001000 : begin
        result = input_776;
      end
      10'b1100001001 : begin
        result = input_777;
      end
      10'b1100001010 : begin
        result = input_778;
      end
      10'b1100001011 : begin
        result = input_779;
      end
      10'b1100001100 : begin
        result = input_780;
      end
      10'b1100001101 : begin
        result = input_781;
      end
      10'b1100001110 : begin
        result = input_782;
      end
      10'b1100001111 : begin
        result = input_783;
      end
      10'b1100010000 : begin
        result = input_784;
      end
      10'b1100010001 : begin
        result = input_785;
      end
      10'b1100010010 : begin
        result = input_786;
      end
      10'b1100010011 : begin
        result = input_787;
      end
      10'b1100010100 : begin
        result = input_788;
      end
      10'b1100010101 : begin
        result = input_789;
      end
      10'b1100010110 : begin
        result = input_790;
      end
      10'b1100010111 : begin
        result = input_791;
      end
      10'b1100011000 : begin
        result = input_792;
      end
      10'b1100011001 : begin
        result = input_793;
      end
      10'b1100011010 : begin
        result = input_794;
      end
      10'b1100011011 : begin
        result = input_795;
      end
      10'b1100011100 : begin
        result = input_796;
      end
      10'b1100011101 : begin
        result = input_797;
      end
      10'b1100011110 : begin
        result = input_798;
      end
      10'b1100011111 : begin
        result = input_799;
      end
      10'b1100100000 : begin
        result = input_800;
      end
      10'b1100100001 : begin
        result = input_801;
      end
      10'b1100100010 : begin
        result = input_802;
      end
      10'b1100100011 : begin
        result = input_803;
      end
      10'b1100100100 : begin
        result = input_804;
      end
      10'b1100100101 : begin
        result = input_805;
      end
      10'b1100100110 : begin
        result = input_806;
      end
      10'b1100100111 : begin
        result = input_807;
      end
      10'b1100101000 : begin
        result = input_808;
      end
      10'b1100101001 : begin
        result = input_809;
      end
      10'b1100101010 : begin
        result = input_810;
      end
      10'b1100101011 : begin
        result = input_811;
      end
      10'b1100101100 : begin
        result = input_812;
      end
      10'b1100101101 : begin
        result = input_813;
      end
      10'b1100101110 : begin
        result = input_814;
      end
      10'b1100101111 : begin
        result = input_815;
      end
      10'b1100110000 : begin
        result = input_816;
      end
      10'b1100110001 : begin
        result = input_817;
      end
      10'b1100110010 : begin
        result = input_818;
      end
      10'b1100110011 : begin
        result = input_819;
      end
      10'b1100110100 : begin
        result = input_820;
      end
      10'b1100110101 : begin
        result = input_821;
      end
      10'b1100110110 : begin
        result = input_822;
      end
      10'b1100110111 : begin
        result = input_823;
      end
      10'b1100111000 : begin
        result = input_824;
      end
      10'b1100111001 : begin
        result = input_825;
      end
      10'b1100111010 : begin
        result = input_826;
      end
      10'b1100111011 : begin
        result = input_827;
      end
      10'b1100111100 : begin
        result = input_828;
      end
      10'b1100111101 : begin
        result = input_829;
      end
      10'b1100111110 : begin
        result = input_830;
      end
      10'b1100111111 : begin
        result = input_831;
      end
      10'b1101000000 : begin
        result = input_832;
      end
      10'b1101000001 : begin
        result = input_833;
      end
      10'b1101000010 : begin
        result = input_834;
      end
      10'b1101000011 : begin
        result = input_835;
      end
      10'b1101000100 : begin
        result = input_836;
      end
      10'b1101000101 : begin
        result = input_837;
      end
      10'b1101000110 : begin
        result = input_838;
      end
      10'b1101000111 : begin
        result = input_839;
      end
      10'b1101001000 : begin
        result = input_840;
      end
      10'b1101001001 : begin
        result = input_841;
      end
      10'b1101001010 : begin
        result = input_842;
      end
      10'b1101001011 : begin
        result = input_843;
      end
      10'b1101001100 : begin
        result = input_844;
      end
      10'b1101001101 : begin
        result = input_845;
      end
      10'b1101001110 : begin
        result = input_846;
      end
      10'b1101001111 : begin
        result = input_847;
      end
      10'b1101010000 : begin
        result = input_848;
      end
      10'b1101010001 : begin
        result = input_849;
      end
      10'b1101010010 : begin
        result = input_850;
      end
      10'b1101010011 : begin
        result = input_851;
      end
      10'b1101010100 : begin
        result = input_852;
      end
      10'b1101010101 : begin
        result = input_853;
      end
      10'b1101010110 : begin
        result = input_854;
      end
      10'b1101010111 : begin
        result = input_855;
      end
      10'b1101011000 : begin
        result = input_856;
      end
      10'b1101011001 : begin
        result = input_857;
      end
      10'b1101011010 : begin
        result = input_858;
      end
      10'b1101011011 : begin
        result = input_859;
      end
      10'b1101011100 : begin
        result = input_860;
      end
      10'b1101011101 : begin
        result = input_861;
      end
      10'b1101011110 : begin
        result = input_862;
      end
      10'b1101011111 : begin
        result = input_863;
      end
      10'b1101100000 : begin
        result = input_864;
      end
      10'b1101100001 : begin
        result = input_865;
      end
      10'b1101100010 : begin
        result = input_866;
      end
      10'b1101100011 : begin
        result = input_867;
      end
      10'b1101100100 : begin
        result = input_868;
      end
      10'b1101100101 : begin
        result = input_869;
      end
      10'b1101100110 : begin
        result = input_870;
      end
      10'b1101100111 : begin
        result = input_871;
      end
      10'b1101101000 : begin
        result = input_872;
      end
      10'b1101101001 : begin
        result = input_873;
      end
      10'b1101101010 : begin
        result = input_874;
      end
      10'b1101101011 : begin
        result = input_875;
      end
      10'b1101101100 : begin
        result = input_876;
      end
      10'b1101101101 : begin
        result = input_877;
      end
      10'b1101101110 : begin
        result = input_878;
      end
      10'b1101101111 : begin
        result = input_879;
      end
      10'b1101110000 : begin
        result = input_880;
      end
      10'b1101110001 : begin
        result = input_881;
      end
      10'b1101110010 : begin
        result = input_882;
      end
      10'b1101110011 : begin
        result = input_883;
      end
      10'b1101110100 : begin
        result = input_884;
      end
      10'b1101110101 : begin
        result = input_885;
      end
      10'b1101110110 : begin
        result = input_886;
      end
      10'b1101110111 : begin
        result = input_887;
      end
      10'b1101111000 : begin
        result = input_888;
      end
      10'b1101111001 : begin
        result = input_889;
      end
      10'b1101111010 : begin
        result = input_890;
      end
      10'b1101111011 : begin
        result = input_891;
      end
      10'b1101111100 : begin
        result = input_892;
      end
      10'b1101111101 : begin
        result = input_893;
      end
      10'b1101111110 : begin
        result = input_894;
      end
      10'b1101111111 : begin
        result = input_895;
      end
      10'b1110000000 : begin
        result = input_896;
      end
      10'b1110000001 : begin
        result = input_897;
      end
      10'b1110000010 : begin
        result = input_898;
      end
      10'b1110000011 : begin
        result = input_899;
      end
      10'b1110000100 : begin
        result = input_900;
      end
      10'b1110000101 : begin
        result = input_901;
      end
      10'b1110000110 : begin
        result = input_902;
      end
      10'b1110000111 : begin
        result = input_903;
      end
      10'b1110001000 : begin
        result = input_904;
      end
      10'b1110001001 : begin
        result = input_905;
      end
      10'b1110001010 : begin
        result = input_906;
      end
      10'b1110001011 : begin
        result = input_907;
      end
      10'b1110001100 : begin
        result = input_908;
      end
      10'b1110001101 : begin
        result = input_909;
      end
      10'b1110001110 : begin
        result = input_910;
      end
      10'b1110001111 : begin
        result = input_911;
      end
      10'b1110010000 : begin
        result = input_912;
      end
      10'b1110010001 : begin
        result = input_913;
      end
      10'b1110010010 : begin
        result = input_914;
      end
      10'b1110010011 : begin
        result = input_915;
      end
      10'b1110010100 : begin
        result = input_916;
      end
      10'b1110010101 : begin
        result = input_917;
      end
      10'b1110010110 : begin
        result = input_918;
      end
      10'b1110010111 : begin
        result = input_919;
      end
      10'b1110011000 : begin
        result = input_920;
      end
      10'b1110011001 : begin
        result = input_921;
      end
      10'b1110011010 : begin
        result = input_922;
      end
      10'b1110011011 : begin
        result = input_923;
      end
      10'b1110011100 : begin
        result = input_924;
      end
      10'b1110011101 : begin
        result = input_925;
      end
      10'b1110011110 : begin
        result = input_926;
      end
      10'b1110011111 : begin
        result = input_927;
      end
      10'b1110100000 : begin
        result = input_928;
      end
      10'b1110100001 : begin
        result = input_929;
      end
      10'b1110100010 : begin
        result = input_930;
      end
      10'b1110100011 : begin
        result = input_931;
      end
      10'b1110100100 : begin
        result = input_932;
      end
      10'b1110100101 : begin
        result = input_933;
      end
      10'b1110100110 : begin
        result = input_934;
      end
      10'b1110100111 : begin
        result = input_935;
      end
      10'b1110101000 : begin
        result = input_936;
      end
      10'b1110101001 : begin
        result = input_937;
      end
      10'b1110101010 : begin
        result = input_938;
      end
      10'b1110101011 : begin
        result = input_939;
      end
      10'b1110101100 : begin
        result = input_940;
      end
      10'b1110101101 : begin
        result = input_941;
      end
      10'b1110101110 : begin
        result = input_942;
      end
      10'b1110101111 : begin
        result = input_943;
      end
      10'b1110110000 : begin
        result = input_944;
      end
      10'b1110110001 : begin
        result = input_945;
      end
      10'b1110110010 : begin
        result = input_946;
      end
      10'b1110110011 : begin
        result = input_947;
      end
      10'b1110110100 : begin
        result = input_948;
      end
      10'b1110110101 : begin
        result = input_949;
      end
      10'b1110110110 : begin
        result = input_950;
      end
      10'b1110110111 : begin
        result = input_951;
      end
      10'b1110111000 : begin
        result = input_952;
      end
      10'b1110111001 : begin
        result = input_953;
      end
      10'b1110111010 : begin
        result = input_954;
      end
      10'b1110111011 : begin
        result = input_955;
      end
      10'b1110111100 : begin
        result = input_956;
      end
      10'b1110111101 : begin
        result = input_957;
      end
      10'b1110111110 : begin
        result = input_958;
      end
      10'b1110111111 : begin
        result = input_959;
      end
      10'b1111000000 : begin
        result = input_960;
      end
      10'b1111000001 : begin
        result = input_961;
      end
      10'b1111000010 : begin
        result = input_962;
      end
      10'b1111000011 : begin
        result = input_963;
      end
      10'b1111000100 : begin
        result = input_964;
      end
      10'b1111000101 : begin
        result = input_965;
      end
      10'b1111000110 : begin
        result = input_966;
      end
      10'b1111000111 : begin
        result = input_967;
      end
      10'b1111001000 : begin
        result = input_968;
      end
      10'b1111001001 : begin
        result = input_969;
      end
      10'b1111001010 : begin
        result = input_970;
      end
      10'b1111001011 : begin
        result = input_971;
      end
      10'b1111001100 : begin
        result = input_972;
      end
      10'b1111001101 : begin
        result = input_973;
      end
      10'b1111001110 : begin
        result = input_974;
      end
      10'b1111001111 : begin
        result = input_975;
      end
      10'b1111010000 : begin
        result = input_976;
      end
      10'b1111010001 : begin
        result = input_977;
      end
      10'b1111010010 : begin
        result = input_978;
      end
      10'b1111010011 : begin
        result = input_979;
      end
      10'b1111010100 : begin
        result = input_980;
      end
      10'b1111010101 : begin
        result = input_981;
      end
      10'b1111010110 : begin
        result = input_982;
      end
      10'b1111010111 : begin
        result = input_983;
      end
      10'b1111011000 : begin
        result = input_984;
      end
      10'b1111011001 : begin
        result = input_985;
      end
      10'b1111011010 : begin
        result = input_986;
      end
      10'b1111011011 : begin
        result = input_987;
      end
      10'b1111011100 : begin
        result = input_988;
      end
      10'b1111011101 : begin
        result = input_989;
      end
      10'b1111011110 : begin
        result = input_990;
      end
      10'b1111011111 : begin
        result = input_991;
      end
      10'b1111100000 : begin
        result = input_992;
      end
      10'b1111100001 : begin
        result = input_993;
      end
      10'b1111100010 : begin
        result = input_994;
      end
      10'b1111100011 : begin
        result = input_995;
      end
      10'b1111100100 : begin
        result = input_996;
      end
      10'b1111100101 : begin
        result = input_997;
      end
      10'b1111100110 : begin
        result = input_998;
      end
      10'b1111100111 : begin
        result = input_999;
      end
      10'b1111101000 : begin
        result = input_1000;
      end
      10'b1111101001 : begin
        result = input_1001;
      end
      10'b1111101010 : begin
        result = input_1002;
      end
      10'b1111101011 : begin
        result = input_1003;
      end
      10'b1111101100 : begin
        result = input_1004;
      end
      10'b1111101101 : begin
        result = input_1005;
      end
      10'b1111101110 : begin
        result = input_1006;
      end
      10'b1111101111 : begin
        result = input_1007;
      end
      10'b1111110000 : begin
        result = input_1008;
      end
      10'b1111110001 : begin
        result = input_1009;
      end
      10'b1111110010 : begin
        result = input_1010;
      end
      10'b1111110011 : begin
        result = input_1011;
      end
      10'b1111110100 : begin
        result = input_1012;
      end
      10'b1111110101 : begin
        result = input_1013;
      end
      10'b1111110110 : begin
        result = input_1014;
      end
      10'b1111110111 : begin
        result = input_1015;
      end
      10'b1111111000 : begin
        result = input_1016;
      end
      10'b1111111001 : begin
        result = input_1017;
      end
      10'b1111111010 : begin
        result = input_1018;
      end
      10'b1111111011 : begin
        result = input_1019;
      end
      10'b1111111100 : begin
        result = input_1020;
      end
      10'b1111111101 : begin
        result = input_1021;
      end
      10'b1111111110 : begin
        result = input_1022;
      end
      default : begin
        result = input_1023;
      end
    endcase
    MUX_s_1_1024_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function automatic [5:0] conv_s2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_s2s_5_6 = {vector[4], vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    nnet_sigmoid_layer4_t_result_t_sigmoid_config5
// ------------------------------------------------------------------


module nnet_sigmoid_layer4_t_result_t_sigmoid_config5 (
  data_rsc_dat, res_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_srst,
      ccs_ccore_en
);
  input [17:0] data_rsc_dat;
  output [17:0] res_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  nnet_sigmoid_layer4_t_result_t_sigmoid_config5_core nnet_sigmoid_layer4_t_result_t_sigmoid_config5_core_inst
      (
      .data_rsc_dat(data_rsc_dat),
      .res_rsc_z(res_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/nnet__dense_large_layer3_t_layer4_t_config4__ca4a50953aa6feccabc41fc32e82972411965_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4a/835166 Production Release
//  HLS Date:       Thu Sep  5 21:35:46 PDT 2019
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Mon Oct 21 13:59:45 2019
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    nnet_dense_large_layer3_t_layer4_t_config4_core
// ------------------------------------------------------------------


module nnet_dense_large_layer3_t_layer4_t_config4_core (
  data_rsc_dat, res_rsc_z, ccs_ccore_clk, ccs_ccore_srst, ccs_ccore_en
);
  input [575:0] data_rsc_dat;
  output [17:0] res_rsc_z;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [575:0] data_rsci_idat;
  reg [17:0] res_rsci_d;
  wire [18:0] nl_res_rsci_d;
  wire [16:0] MultLoop_acc_97_itm_23_7;
  wire [17:0] MultLoop_acc_141_itm_18_1;

  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_30_nl;
  wire[21:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_30_nl;
  wire[17:0] MultLoop_acc_128_nl;
  wire[18:0] nl_MultLoop_acc_128_nl;
  wire[22:0] MultLoop_acc_85_nl;
  wire[24:0] nl_MultLoop_acc_85_nl;
  wire[17:0] MultLoop_acc_83_nl;
  wire[18:0] nl_MultLoop_acc_83_nl;
  wire[9:0] MultLoop_acc_127_nl;
  wire[10:0] nl_MultLoop_acc_127_nl;
  wire[18:0] MultLoop_acc_130_nl;
  wire[19:0] nl_MultLoop_acc_130_nl;
  wire[18:0] MultLoop_acc_129_nl;
  wire[19:0] nl_MultLoop_acc_129_nl;
  wire[20:0] MultLoop_acc_86_nl;
  wire[21:0] nl_MultLoop_acc_86_nl;
  wire[17:0] MultLoop_acc_132_nl;
  wire[18:0] nl_MultLoop_acc_132_nl;
  wire[18:0] MultLoop_acc_131_nl;
  wire[19:0] nl_MultLoop_acc_131_nl;
  wire[22:0] MultLoop_acc_89_nl;
  wire[24:0] nl_MultLoop_acc_89_nl;
  wire[20:0] MultLoop_acc_135_nl;
  wire[21:0] nl_MultLoop_acc_135_nl;
  wire[17:0] MultLoop_acc_134_nl;
  wire[18:0] nl_MultLoop_acc_134_nl;
  wire[20:0] MultLoop_acc_92_nl;
  wire[21:0] nl_MultLoop_acc_92_nl;
  wire[9:0] MultLoop_acc_133_nl;
  wire[10:0] nl_MultLoop_acc_133_nl;
  wire[16:0] MultLoop_acc_137_nl;
  wire[17:0] nl_MultLoop_acc_137_nl;
  wire[18:0] MultLoop_acc_138_nl;
  wire[19:0] nl_MultLoop_acc_138_nl;
  wire[22:0] MultLoop_acc_99_nl;
  wire[24:0] nl_MultLoop_acc_99_nl;
  wire[17:0] MultLoop_acc_139_nl;
  wire[18:0] nl_MultLoop_acc_139_nl;
  wire[22:0] MultLoop_acc_102_nl;
  wire[23:0] nl_MultLoop_acc_102_nl;
  wire[19:0] MultLoop_acc_101_nl;
  wire[21:0] nl_MultLoop_acc_101_nl;
  wire[16:0] MultLoop_acc_142_nl;
  wire[17:0] nl_MultLoop_acc_142_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_9_nl;
  wire[18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_9_nl;
  wire[27:0] MultLoop_acc_34_nl;
  wire[29:0] nl_MultLoop_acc_34_nl;
  wire[9:0] MultLoop_acc_149_nl;
  wire[10:0] nl_MultLoop_acc_149_nl;
  wire[21:0] MultLoop_acc_45_nl;
  wire[22:0] nl_MultLoop_acc_45_nl;
  wire[19:0] MultLoop_acc_126_nl;
  wire[21:0] nl_MultLoop_acc_126_nl;
  wire[19:0] MultLoop_acc_148_nl;
  wire[20:0] nl_MultLoop_acc_148_nl;
  wire[17:0] MultLoop_acc_147_nl;
  wire[18:0] nl_MultLoop_acc_147_nl;
  wire[20:0] MultLoop_acc_119_nl;
  wire[21:0] nl_MultLoop_acc_119_nl;
  wire[22:0] MultLoop_acc_44_nl;
  wire[23:0] nl_MultLoop_acc_44_nl;
  wire[19:0] MultLoop_acc_122_nl;
  wire[21:0] nl_MultLoop_acc_122_nl;
  wire[21:0] MultLoop_acc_41_nl;
  wire[22:0] nl_MultLoop_acc_41_nl;
  wire[19:0] MultLoop_acc_109_nl;
  wire[20:0] nl_MultLoop_acc_109_nl;
  wire[17:0] MultLoop_acc_108_nl;
  wire[18:0] nl_MultLoop_acc_108_nl;
  wire[25:0] MultLoop_acc_42_nl;
  wire[26:0] nl_MultLoop_acc_42_nl;
  wire[22:0] MultLoop_acc_112_nl;
  wire[24:0] nl_MultLoop_acc_112_nl;
  wire[9:0] MultLoop_acc_143_nl;
  wire[10:0] nl_MultLoop_acc_143_nl;
  wire[22:0] MultLoop_acc_43_nl;
  wire[23:0] nl_MultLoop_acc_43_nl;
  wire[19:0] MultLoop_acc_115_nl;
  wire[21:0] nl_MultLoop_acc_115_nl;
  wire[10:0] MultLoop_acc_144_nl;
  wire[11:0] nl_MultLoop_acc_144_nl;
  wire[17:0] MultLoop_acc_146_nl;
  wire[18:0] nl_MultLoop_acc_146_nl;
  wire[23:0] MultLoop_acc_118_nl;
  wire[24:0] nl_MultLoop_acc_118_nl;
  wire[20:0] MultLoop_acc_117_nl;
  wire[21:0] nl_MultLoop_acc_117_nl;
  wire[8:0] MultLoop_acc_145_nl;
  wire[9:0] nl_MultLoop_acc_145_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_nl;
  wire[19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_25_nl;
  wire[18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_25_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_18_nl;
  wire[19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_18_nl;
  wire[17:0] MultLoop_acc_157_nl;
  wire[18:0] nl_MultLoop_acc_157_nl;
  wire[19:0] MultLoop_acc_64_nl;
  wire[20:0] nl_MultLoop_acc_64_nl;
  wire[17:0] MultLoop_acc_63_nl;
  wire[18:0] nl_MultLoop_acc_63_nl;
  wire[9:0] MultLoop_acc_156_nl;
  wire[10:0] nl_MultLoop_acc_156_nl;
  wire[17:0] MultLoop_acc_159_nl;
  wire[18:0] nl_MultLoop_acc_159_nl;
  wire[21:0] MultLoop_acc_68_nl;
  wire[22:0] nl_MultLoop_acc_68_nl;
  wire[19:0] MultLoop_acc_67_nl;
  wire[21:0] nl_MultLoop_acc_67_nl;
  wire[9:0] MultLoop_acc_158_nl;
  wire[10:0] nl_MultLoop_acc_158_nl;
  wire[17:0] MultLoop_acc_161_nl;
  wire[18:0] nl_MultLoop_acc_161_nl;
  wire[24:0] MultLoop_acc_72_nl;
  wire[25:0] nl_MultLoop_acc_72_nl;
  wire[21:0] MultLoop_acc_71_nl;
  wire[23:0] nl_MultLoop_acc_71_nl;
  wire[9:0] MultLoop_acc_160_nl;
  wire[10:0] nl_MultLoop_acc_160_nl;
  wire[19:0] MultLoop_acc_163_nl;
  wire[20:0] nl_MultLoop_acc_163_nl;
  wire[17:0] MultLoop_acc_162_nl;
  wire[18:0] nl_MultLoop_acc_162_nl;
  wire[22:0] MultLoop_acc_74_nl;
  wire[23:0] nl_MultLoop_acc_74_nl;
  wire[19:0] MultLoop_acc_73_nl;
  wire[20:0] nl_MultLoop_acc_73_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_17_nl;
  wire[18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_17_nl;
  wire[24:0] MultLoop_acc_38_nl;
  wire[25:0] nl_MultLoop_acc_38_nl;
  wire[22:0] MultLoop_acc_78_nl;
  wire[23:0] nl_MultLoop_acc_78_nl;
  wire[17:0] MultLoop_acc_77_nl;
  wire[18:0] nl_MultLoop_acc_77_nl;
  wire[9:0] MultLoop_acc_164_nl;
  wire[10:0] nl_MultLoop_acc_164_nl;
  wire[24:0] MultLoop_acc_39_nl;
  wire[25:0] nl_MultLoop_acc_39_nl;
  wire[21:0] MultLoop_acc_81_nl;
  wire[23:0] nl_MultLoop_acc_81_nl;
  wire[10:0] MultLoop_acc_165_nl;
  wire[11:0] nl_MultLoop_acc_165_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_26_nl;
  wire[20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_26_nl;
  wire[18:0] MultLoop_acc_152_nl;
  wire[19:0] nl_MultLoop_acc_152_nl;
  wire[22:0] MultLoop_acc_51_nl;
  wire[23:0] nl_MultLoop_acc_51_nl;
  wire[24:0] MultLoop_acc_21_nl;
  wire[25:0] nl_MultLoop_acc_21_nl;
  wire[21:0] MultLoop_acc_53_nl;
  wire[23:0] nl_MultLoop_acc_53_nl;
  wire[15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_2_nl;
  wire[16:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_2_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_nor_nl;
  wire[20:0] MultLoop_acc_nl;
  wire[21:0] nl_MultLoop_acc_nl;
  wire[17:0] MultLoop_acc_47_nl;
  wire[18:0] nl_MultLoop_acc_47_nl;
  wire[12:0] MultLoop_acc_150_nl;
  wire[13:0] nl_MultLoop_acc_150_nl;
  wire[17:0] MultLoop_acc_14_nl;
  wire[18:0] nl_MultLoop_acc_14_nl;
  wire[21:0] MultLoop_acc_35_nl;
  wire[22:0] nl_MultLoop_acc_35_nl;
  wire[19:0] MultLoop_acc_50_nl;
  wire[20:0] nl_MultLoop_acc_50_nl;
  wire[17:0] MultLoop_acc_49_nl;
  wire[18:0] nl_MultLoop_acc_49_nl;
  wire[11:0] MultLoop_acc_151_nl;
  wire[12:0] nl_MultLoop_acc_151_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_19_nl;
  wire[19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_19_nl;
  wire[25:0] MultLoop_acc_22_nl;
  wire[26:0] nl_MultLoop_acc_22_nl;
  wire[20:0] MultLoop_acc_54_nl;
  wire[21:0] nl_MultLoop_acc_54_nl;
  wire[21:0] MultLoop_acc_37_nl;
  wire[22:0] nl_MultLoop_acc_37_nl;
  wire[17:0] MultLoop_acc_56_nl;
  wire[18:0] nl_MultLoop_acc_56_nl;
  wire[12:0] MultLoop_acc_153_nl;
  wire[13:0] nl_MultLoop_acc_153_nl;
  wire[25:0] MultLoop_acc_26_nl;
  wire[26:0] nl_MultLoop_acc_26_nl;
  wire[24:0] MultLoop_acc_58_nl;
  wire[26:0] nl_MultLoop_acc_58_nl;
  wire[17:0] MultLoop_acc_155_nl;
  wire[18:0] nl_MultLoop_acc_155_nl;
  wire[23:0] MultLoop_acc_61_nl;
  wire[24:0] nl_MultLoop_acc_61_nl;
  wire[19:0] MultLoop_acc_60_nl;
  wire[20:0] nl_MultLoop_acc_60_nl;
  wire[10:0] MultLoop_acc_154_nl;
  wire[11:0] nl_MultLoop_acc_154_nl;
  wire[23:0] MultLoop_acc_97_nl;
  wire[25:0] nl_MultLoop_acc_97_nl;
  wire[17:0] MultLoop_acc_95_nl;
  wire[18:0] nl_MultLoop_acc_95_nl;
  wire[7:0] MultLoop_acc_136_nl;
  wire[8:0] nl_MultLoop_acc_136_nl;
  wire[18:0] MultLoop_acc_141_nl;
  wire[19:0] nl_MultLoop_acc_141_nl;
  wire[23:0] MultLoop_acc_106_nl;
  wire[25:0] nl_MultLoop_acc_106_nl;
  wire[7:0] MultLoop_acc_140_nl;
  wire[8:0] nl_MultLoop_acc_140_nl;

  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd8),
  .width(32'sd576)) data_rsci (
      .dat(data_rsc_dat),
      .idat(data_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd9),
  .width(32'sd18)) res_rsci (
      .d(res_rsci_d),
      .z(res_rsc_z)
    );
  assign nl_MultLoop_acc_136_nl = conv_s2s_7_8(data_rsci_idat[179:173]) + 8'b00000001;
  assign MultLoop_acc_136_nl = nl_MultLoop_acc_136_nl[7:0];
  assign nl_MultLoop_acc_95_nl = (~ (data_rsci_idat[179:162])) + conv_s2s_16_18({(MultLoop_acc_136_nl)
      , (data_rsci_idat[172:165])});
  assign MultLoop_acc_95_nl = nl_MultLoop_acc_95_nl[17:0];
  assign nl_MultLoop_acc_97_nl = ({(data_rsci_idat[179:162]) , 6'b010000}) + conv_s2s_22_24({(~
      (data_rsci_idat[179:162])) , 4'b0001}) + conv_s2s_18_24(MultLoop_acc_95_nl);
  assign MultLoop_acc_97_nl = nl_MultLoop_acc_97_nl[23:0];
  assign MultLoop_acc_97_itm_23_7 = readslicef_24_17_7((MultLoop_acc_97_nl));
  assign nl_MultLoop_acc_140_nl = conv_s2s_7_8(data_rsci_idat[233:227]) + 8'b00000001;
  assign MultLoop_acc_140_nl = nl_MultLoop_acc_140_nl[7:0];
  assign nl_MultLoop_acc_106_nl = conv_s2s_23_24({(data_rsci_idat[233:216]) , 5'b00000})
      + conv_s2s_21_24({(data_rsci_idat[233:216]) , 3'b000}) + conv_s2s_18_24(data_rsci_idat[233:216])
      + conv_s2s_17_24({(MultLoop_acc_140_nl) , (data_rsci_idat[226:218])});
  assign MultLoop_acc_106_nl = nl_MultLoop_acc_106_nl[23:0];
  assign nl_MultLoop_acc_141_nl = conv_s2u_18_19(data_rsci_idat[233:216]) + conv_s2u_17_19(readslicef_24_17_7((MultLoop_acc_106_nl)));
  assign MultLoop_acc_141_nl = nl_MultLoop_acc_141_nl[18:0];
  assign MultLoop_acc_141_itm_18_1 = readslicef_19_18_1((MultLoop_acc_141_nl));
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      res_rsci_d <= 18'b000000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      res_rsci_d <= nl_res_rsci_d[17:0];
    end
  end
  assign nl_MultLoop_acc_127_nl = conv_s2s_9_10(data_rsci_idat[53:45]) + 10'b0000000001;
  assign MultLoop_acc_127_nl = nl_MultLoop_acc_127_nl[9:0];
  assign nl_MultLoop_acc_83_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_17_18({(MultLoop_acc_127_nl)
      , (data_rsci_idat[44:38])});
  assign MultLoop_acc_83_nl = nl_MultLoop_acc_83_nl[17:0];
  assign nl_MultLoop_acc_85_nl = ({(data_rsci_idat[53:36]) , 5'b01000}) + conv_s2s_21_23({(~
      (data_rsci_idat[53:36])) , 3'b001}) + conv_s2s_18_23(MultLoop_acc_83_nl);
  assign MultLoop_acc_85_nl = nl_MultLoop_acc_85_nl[22:0];
  assign nl_MultLoop_acc_128_nl = conv_s2u_16_18(readslicef_23_16_7((MultLoop_acc_85_nl)))
      + (~ (data_rsci_idat[53:36]));
  assign MultLoop_acc_128_nl = nl_MultLoop_acc_128_nl[17:0];
  assign nl_MultLoop_acc_86_nl = ({(data_rsci_idat[107:90]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[107:90]));
  assign MultLoop_acc_86_nl = nl_MultLoop_acc_86_nl[20:0];
  assign nl_MultLoop_acc_129_nl = conv_s2u_18_19(data_rsci_idat[107:90]) + conv_s2u_14_19(readslicef_21_14_7((MultLoop_acc_86_nl)));
  assign MultLoop_acc_129_nl = nl_MultLoop_acc_129_nl[18:0];
  assign nl_MultLoop_acc_130_nl = conv_s2u_17_19(readslicef_19_17_2((MultLoop_acc_129_nl)))
      + conv_s2u_18_19(data_rsci_idat[107:90]);
  assign MultLoop_acc_130_nl = nl_MultLoop_acc_130_nl[18:0];
  assign nl_MultLoop_acc_89_nl = ({(data_rsci_idat[125:108]) , 5'b01000}) + conv_s2s_21_23({(~
      (data_rsci_idat[125:108])) , 3'b001}) + conv_s2s_18_23(~ (data_rsci_idat[125:108]));
  assign MultLoop_acc_89_nl = nl_MultLoop_acc_89_nl[22:0];
  assign nl_MultLoop_acc_131_nl = conv_s2u_18_19(data_rsci_idat[125:108]) + conv_s2u_16_19(readslicef_23_16_7((MultLoop_acc_89_nl)));
  assign MultLoop_acc_131_nl = nl_MultLoop_acc_131_nl[18:0];
  assign nl_MultLoop_acc_132_nl = conv_s2u_17_18(readslicef_19_17_2((MultLoop_acc_131_nl)))
      + (data_rsci_idat[125:108]);
  assign MultLoop_acc_132_nl = nl_MultLoop_acc_132_nl[17:0];
  assign nl_MultLoop_acc_133_nl =  -conv_s2s_9_10(data_rsci_idat[143:135]);
  assign MultLoop_acc_133_nl = nl_MultLoop_acc_133_nl[9:0];
  assign nl_MultLoop_acc_92_nl = ({(data_rsci_idat[143:126]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_133_nl)
      , (~ (data_rsci_idat[134:126]))});
  assign MultLoop_acc_92_nl = nl_MultLoop_acc_92_nl[20:0];
  assign nl_MultLoop_acc_134_nl = (~ (data_rsci_idat[143:126])) + conv_s2s_14_18(readslicef_21_14_7((MultLoop_acc_92_nl)));
  assign MultLoop_acc_134_nl = nl_MultLoop_acc_134_nl[17:0];
  assign nl_MultLoop_acc_135_nl = conv_s2u_18_21(MultLoop_acc_134_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[143:126])) , 2'b01});
  assign MultLoop_acc_135_nl = nl_MultLoop_acc_135_nl[20:0];
  assign nl_MultLoop_acc_137_nl = conv_s2u_16_17(MultLoop_acc_97_itm_23_7[16:1])
      + (~ (data_rsci_idat[178:162]));
  assign MultLoop_acc_137_nl = nl_MultLoop_acc_137_nl[16:0];
  assign nl_MultLoop_acc_99_nl = ({(data_rsci_idat[197:180]) , 5'b00100}) + conv_s2s_20_23({(~
      (data_rsci_idat[197:180])) , 2'b01}) + conv_s2s_18_23(~ (data_rsci_idat[197:180]));
  assign MultLoop_acc_99_nl = nl_MultLoop_acc_99_nl[22:0];
  assign nl_MultLoop_acc_138_nl = conv_s2u_15_19(readslicef_23_15_8((MultLoop_acc_99_nl)))
      + conv_s2u_18_19(data_rsci_idat[197:180]);
  assign MultLoop_acc_138_nl = nl_MultLoop_acc_138_nl[18:0];
  assign nl_MultLoop_acc_101_nl = ({(~ (data_rsci_idat[215:198])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[215:198])
      + conv_s2s_15_20(data_rsci_idat[215:201]);
  assign MultLoop_acc_101_nl = nl_MultLoop_acc_101_nl[19:0];
  assign nl_MultLoop_acc_102_nl = ({(data_rsci_idat[215:198]) , 5'b00100}) + conv_s2s_20_23(MultLoop_acc_101_nl);
  assign MultLoop_acc_102_nl = nl_MultLoop_acc_102_nl[22:0];
  assign nl_MultLoop_acc_139_nl = conv_s2u_16_18(readslicef_23_16_7((MultLoop_acc_102_nl)))
      + (data_rsci_idat[215:198]);
  assign MultLoop_acc_139_nl = nl_MultLoop_acc_139_nl[17:0];
  assign nl_MultLoop_acc_142_nl = (MultLoop_acc_141_itm_18_1[17:1]) + (~ (data_rsci_idat[232:216]));
  assign MultLoop_acc_142_nl = nl_MultLoop_acc_142_nl[16:0];
  assign nl_MultLoop_acc_149_nl =  -conv_s2s_9_10(data_rsci_idat[539:531]);
  assign MultLoop_acc_149_nl = nl_MultLoop_acc_149_nl[9:0];
  assign nl_MultLoop_acc_34_nl = conv_s2s_27_28({(~ (data_rsci_idat[539:522])) ,
      9'b001000000}) + conv_s2s_24_28({(~ (data_rsci_idat[539:522])) , 6'b000001})
      + conv_s2s_19_28({(MultLoop_acc_149_nl) , (~ (data_rsci_idat[530:522]))});
  assign MultLoop_acc_34_nl = nl_MultLoop_acc_34_nl[27:0];
  assign nl_MultLoop_acc_126_nl = ({(~ (data_rsci_idat[575:558])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[575:558])
      + conv_s2s_15_20(data_rsci_idat[575:561]);
  assign MultLoop_acc_126_nl = nl_MultLoop_acc_126_nl[19:0];
  assign nl_MultLoop_acc_45_nl = conv_s2u_20_22(MultLoop_acc_126_nl) + ({(data_rsci_idat[575:558])
      , 4'b0100});
  assign MultLoop_acc_45_nl = nl_MultLoop_acc_45_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_9_nl = (readslicef_28_18_10((MultLoop_acc_34_nl)))
      + (readslicef_22_18_4((MultLoop_acc_45_nl)));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_9_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_9_nl[17:0];
  assign nl_MultLoop_acc_119_nl = ({(data_rsci_idat[485:468]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[485:468]));
  assign MultLoop_acc_119_nl = nl_MultLoop_acc_119_nl[20:0];
  assign nl_MultLoop_acc_147_nl = (~ (data_rsci_idat[485:468])) + conv_s2s_13_18(readslicef_21_13_8((MultLoop_acc_119_nl)));
  assign MultLoop_acc_147_nl = nl_MultLoop_acc_147_nl[17:0];
  assign nl_MultLoop_acc_148_nl = conv_s2u_18_20(MultLoop_acc_147_nl) + ({(data_rsci_idat[485:468])
      , 2'b01});
  assign MultLoop_acc_148_nl = nl_MultLoop_acc_148_nl[19:0];
  assign nl_MultLoop_acc_122_nl = ({(~ (data_rsci_idat[521:504])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[521:504])
      + conv_s2s_15_20(data_rsci_idat[521:507]);
  assign MultLoop_acc_122_nl = nl_MultLoop_acc_122_nl[19:0];
  assign nl_MultLoop_acc_44_nl = conv_s2u_20_23(MultLoop_acc_122_nl) + ({(data_rsci_idat[521:504])
      , 5'b00100});
  assign MultLoop_acc_44_nl = nl_MultLoop_acc_44_nl[22:0];
  assign nl_MultLoop_acc_108_nl = (~ (data_rsci_idat[251:234])) + conv_s2s_15_18(data_rsci_idat[251:237]);
  assign MultLoop_acc_108_nl = nl_MultLoop_acc_108_nl[17:0];
  assign nl_MultLoop_acc_109_nl = ({(data_rsci_idat[251:234]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_108_nl);
  assign MultLoop_acc_109_nl = nl_MultLoop_acc_109_nl[19:0];
  assign nl_MultLoop_acc_41_nl = conv_s2u_20_22(MultLoop_acc_109_nl) + ({(data_rsci_idat[251:234])
      , 4'b0000});
  assign MultLoop_acc_41_nl = nl_MultLoop_acc_41_nl[21:0];
  assign nl_MultLoop_acc_143_nl = conv_s2s_9_10(data_rsci_idat[269:261]) + 10'b0000000001;
  assign MultLoop_acc_143_nl = nl_MultLoop_acc_143_nl[9:0];
  assign nl_MultLoop_acc_112_nl = ({(~ (data_rsci_idat[269:252])) , 5'b00000}) +
      conv_s2s_18_23(data_rsci_idat[269:252]) + conv_s2s_17_23({(MultLoop_acc_143_nl)
      , (data_rsci_idat[260:254])});
  assign MultLoop_acc_112_nl = nl_MultLoop_acc_112_nl[22:0];
  assign nl_MultLoop_acc_42_nl = conv_s2u_23_26(MultLoop_acc_112_nl) + conv_s2u_25_26({(~
      (data_rsci_idat[269:252])) , 7'b0100000});
  assign MultLoop_acc_42_nl = nl_MultLoop_acc_42_nl[25:0];
  assign nl_MultLoop_acc_144_nl = conv_s2s_10_11(data_rsci_idat[323:314]) + 11'b00000000001;
  assign MultLoop_acc_144_nl = nl_MultLoop_acc_144_nl[10:0];
  assign nl_MultLoop_acc_115_nl = ({(~ (data_rsci_idat[323:306])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[323:306])
      + conv_s2s_15_20({(MultLoop_acc_144_nl) , (data_rsci_idat[313:310])});
  assign MultLoop_acc_115_nl = nl_MultLoop_acc_115_nl[19:0];
  assign nl_MultLoop_acc_43_nl = conv_s2u_20_23(MultLoop_acc_115_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[323:306])) , 4'b0100});
  assign MultLoop_acc_43_nl = nl_MultLoop_acc_43_nl[22:0];
  assign nl_MultLoop_acc_145_nl =  -conv_s2s_8_9(data_rsci_idat[341:334]);
  assign MultLoop_acc_145_nl = nl_MultLoop_acc_145_nl[8:0];
  assign nl_MultLoop_acc_117_nl = ({(data_rsci_idat[341:324]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_145_nl)
      , (~ (data_rsci_idat[333:324]))});
  assign MultLoop_acc_117_nl = nl_MultLoop_acc_117_nl[20:0];
  assign nl_MultLoop_acc_118_nl = conv_s2s_23_24({(data_rsci_idat[341:324]) , 5'b00000})
      + conv_s2s_21_24(MultLoop_acc_117_nl);
  assign MultLoop_acc_118_nl = nl_MultLoop_acc_118_nl[23:0];
  assign nl_MultLoop_acc_146_nl = conv_s2u_14_18(readslicef_24_14_10((MultLoop_acc_118_nl)))
      + (~ (data_rsci_idat[341:324]));
  assign MultLoop_acc_146_nl = nl_MultLoop_acc_146_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_30_nl = (MultLoop_acc_128_nl)
      + (readslicef_19_18_1((MultLoop_acc_130_nl))) + (MultLoop_acc_132_nl) + (readslicef_21_18_3((MultLoop_acc_135_nl)))
      + ({(MultLoop_acc_137_nl) , (MultLoop_acc_97_itm_23_7[0])}) + (readslicef_19_18_1((MultLoop_acc_138_nl)))
      + (MultLoop_acc_139_nl) + ({(MultLoop_acc_142_nl) , (MultLoop_acc_141_itm_18_1[0])})
      + (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_9_nl) + (readslicef_20_18_2((MultLoop_acc_148_nl)))
      + (readslicef_23_18_5((MultLoop_acc_44_nl))) + (readslicef_22_18_4((MultLoop_acc_41_nl)))
      + (readslicef_26_18_8((MultLoop_acc_42_nl))) + (readslicef_23_18_5((MultLoop_acc_43_nl)))
      + (MultLoop_acc_146_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_30_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_30_nl[17:0];
  assign nl_MultLoop_acc_156_nl = conv_s2s_9_10(data_rsci_idat[431:423]) + 10'b0000000001;
  assign MultLoop_acc_156_nl = nl_MultLoop_acc_156_nl[9:0];
  assign nl_MultLoop_acc_63_nl = (~ (data_rsci_idat[431:414])) + conv_s2s_17_18({(MultLoop_acc_156_nl)
      , (data_rsci_idat[422:416])});
  assign MultLoop_acc_63_nl = nl_MultLoop_acc_63_nl[17:0];
  assign nl_MultLoop_acc_64_nl = ({(data_rsci_idat[431:414]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_63_nl);
  assign MultLoop_acc_64_nl = nl_MultLoop_acc_64_nl[19:0];
  assign nl_MultLoop_acc_157_nl = conv_s2u_13_18(readslicef_20_13_7((MultLoop_acc_64_nl)))
      + (~ (data_rsci_idat[431:414]));
  assign MultLoop_acc_157_nl = nl_MultLoop_acc_157_nl[17:0];
  assign nl_MultLoop_acc_158_nl = conv_s2s_9_10(data_rsci_idat[449:441]) + 10'b0000000001;
  assign MultLoop_acc_158_nl = nl_MultLoop_acc_158_nl[9:0];
  assign nl_MultLoop_acc_67_nl = ({(~ (data_rsci_idat[449:432])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[449:432])
      + conv_s2s_16_20({(MultLoop_acc_158_nl) , (data_rsci_idat[440:435])});
  assign MultLoop_acc_67_nl = nl_MultLoop_acc_67_nl[19:0];
  assign nl_MultLoop_acc_68_nl = ({(data_rsci_idat[449:432]) , 4'b0100}) + conv_s2s_20_22(MultLoop_acc_67_nl);
  assign MultLoop_acc_68_nl = nl_MultLoop_acc_68_nl[21:0];
  assign nl_MultLoop_acc_159_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_68_nl)))
      + (~ (data_rsci_idat[449:432]));
  assign MultLoop_acc_159_nl = nl_MultLoop_acc_159_nl[17:0];
  assign nl_MultLoop_acc_160_nl =  -conv_s2s_9_10(data_rsci_idat[467:459]);
  assign MultLoop_acc_160_nl = nl_MultLoop_acc_160_nl[9:0];
  assign nl_MultLoop_acc_71_nl = ({(data_rsci_idat[467:450]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[467:450])) , 2'b01}) + conv_s2s_19_22({(MultLoop_acc_160_nl)
      , (~ (data_rsci_idat[458:450]))});
  assign MultLoop_acc_71_nl = nl_MultLoop_acc_71_nl[21:0];
  assign nl_MultLoop_acc_72_nl = conv_s2s_24_25({(data_rsci_idat[467:450]) , 6'b000000})
      + conv_s2s_22_25(MultLoop_acc_71_nl);
  assign MultLoop_acc_72_nl = nl_MultLoop_acc_72_nl[24:0];
  assign nl_MultLoop_acc_161_nl = conv_s2u_16_18(readslicef_25_16_9((MultLoop_acc_72_nl)))
      + (~ (data_rsci_idat[467:450]));
  assign MultLoop_acc_161_nl = nl_MultLoop_acc_161_nl[17:0];
  assign nl_MultLoop_acc_73_nl = ({(data_rsci_idat[503:486]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[503:486]));
  assign MultLoop_acc_73_nl = nl_MultLoop_acc_73_nl[19:0];
  assign nl_MultLoop_acc_74_nl = conv_s2s_22_23({(data_rsci_idat[503:486]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_73_nl);
  assign MultLoop_acc_74_nl = nl_MultLoop_acc_74_nl[22:0];
  assign nl_MultLoop_acc_162_nl = (~ (data_rsci_idat[503:486])) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_74_nl)));
  assign MultLoop_acc_162_nl = nl_MultLoop_acc_162_nl[17:0];
  assign nl_MultLoop_acc_163_nl = conv_s2u_18_20(MultLoop_acc_162_nl) + ({(data_rsci_idat[503:486])
      , 2'b01});
  assign MultLoop_acc_163_nl = nl_MultLoop_acc_163_nl[19:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_18_nl = conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_157_nl)))
      + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_159_nl))) + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_161_nl)))
      + conv_s2s_17_18(readslicef_20_17_3((MultLoop_acc_163_nl)));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_18_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_18_nl[17:0];
  assign nl_MultLoop_acc_164_nl = conv_s2s_9_10(data_rsci_idat[17:9]) + 10'b0000000001;
  assign MultLoop_acc_164_nl = nl_MultLoop_acc_164_nl[9:0];
  assign nl_MultLoop_acc_77_nl = (~ (data_rsci_idat[17:0])) + conv_s2s_17_18({(MultLoop_acc_164_nl)
      , (data_rsci_idat[8:2])});
  assign MultLoop_acc_77_nl = nl_MultLoop_acc_77_nl[17:0];
  assign nl_MultLoop_acc_78_nl = conv_s2s_22_23({(~ (data_rsci_idat[17:0])) , 4'b0001})
      + conv_s2s_18_23(MultLoop_acc_77_nl);
  assign MultLoop_acc_78_nl = nl_MultLoop_acc_78_nl[22:0];
  assign nl_MultLoop_acc_38_nl = conv_s2u_23_25(MultLoop_acc_78_nl) + ({(~ (data_rsci_idat[17:0]))
      , 7'b0010000});
  assign MultLoop_acc_38_nl = nl_MultLoop_acc_38_nl[24:0];
  assign nl_MultLoop_acc_165_nl = conv_s2s_10_11(data_rsci_idat[35:26]) + 11'b00000000001;
  assign MultLoop_acc_165_nl = nl_MultLoop_acc_165_nl[10:0];
  assign nl_MultLoop_acc_81_nl = ({(~ (data_rsci_idat[35:18])) , 4'b0000}) + conv_s2s_18_22(data_rsci_idat[35:18])
      + conv_s2s_17_22({(MultLoop_acc_165_nl) , (data_rsci_idat[25:20])});
  assign MultLoop_acc_81_nl = nl_MultLoop_acc_81_nl[21:0];
  assign nl_MultLoop_acc_39_nl = conv_s2u_22_25(MultLoop_acc_81_nl) + conv_s2u_24_25({(~
      (data_rsci_idat[35:18])) , 6'b010000});
  assign MultLoop_acc_39_nl = nl_MultLoop_acc_39_nl[24:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_17_nl = (readslicef_25_18_7((MultLoop_acc_38_nl)))
      + (readslicef_25_18_7((MultLoop_acc_39_nl)));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_17_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_17_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_25_nl = (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_18_nl)
      + (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_17_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_25_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_25_nl[17:0];
  assign nl_MultLoop_acc_51_nl = ({(data_rsci_idat[89:72]) , 5'b00001}) + conv_s2s_18_23(~
      (data_rsci_idat[89:72]));
  assign MultLoop_acc_51_nl = nl_MultLoop_acc_51_nl[22:0];
  assign nl_MultLoop_acc_152_nl = conv_s2u_15_19(readslicef_23_15_8((MultLoop_acc_51_nl)))
      + conv_s2u_18_19(data_rsci_idat[89:72]);
  assign MultLoop_acc_152_nl = nl_MultLoop_acc_152_nl[18:0];
  assign nl_MultLoop_acc_53_nl = ({(data_rsci_idat[287:270]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[287:270])) , 2'b01}) + conv_s2s_18_22(~ (data_rsci_idat[287:270]));
  assign MultLoop_acc_53_nl = nl_MultLoop_acc_53_nl[21:0];
  assign nl_MultLoop_acc_21_nl = conv_s2s_22_25(MultLoop_acc_53_nl) + conv_s2s_24_25({(data_rsci_idat[287:270])
      , 6'b000000});
  assign MultLoop_acc_21_nl = nl_MultLoop_acc_21_nl[24:0];
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_nor_nl = ~((data_rsci_idat[398:396]!=3'b000));
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_2_nl = conv_s2s_15_16(~
      (data_rsci_idat[413:399])) + conv_u2s_7_16({6'b110010 , (nnet_product_input_t_config2_weight_t_config2_accum_t_nor_nl)});
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_2_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_2_nl[15:0];
  assign nl_MultLoop_acc_150_nl = conv_s2s_12_13(data_rsci_idat[71:60]) + 13'b0000000000001;
  assign MultLoop_acc_150_nl = nl_MultLoop_acc_150_nl[12:0];
  assign nl_MultLoop_acc_47_nl = (~ (data_rsci_idat[71:54])) + conv_s2s_15_18({(MultLoop_acc_150_nl)
      , (data_rsci_idat[59:58])});
  assign MultLoop_acc_47_nl = nl_MultLoop_acc_47_nl[17:0];
  assign nl_MultLoop_acc_nl = conv_s2u_18_21(MultLoop_acc_47_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[71:54])) , 2'b01});
  assign MultLoop_acc_nl = nl_MultLoop_acc_nl[20:0];
  assign nl_MultLoop_acc_14_nl = conv_s2u_15_18(data_rsci_idat[161:147]) - (data_rsci_idat[161:144]);
  assign MultLoop_acc_14_nl = nl_MultLoop_acc_14_nl[17:0];
  assign nl_MultLoop_acc_151_nl = conv_s2s_11_12(data_rsci_idat[557:547]) + 12'b000000000001;
  assign MultLoop_acc_151_nl = nl_MultLoop_acc_151_nl[11:0];
  assign nl_MultLoop_acc_49_nl = (~ (data_rsci_idat[557:540])) + conv_s2s_16_18({(MultLoop_acc_151_nl)
      , (data_rsci_idat[546:543])});
  assign MultLoop_acc_49_nl = nl_MultLoop_acc_49_nl[17:0];
  assign nl_MultLoop_acc_50_nl = ({(data_rsci_idat[557:540]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_49_nl);
  assign MultLoop_acc_50_nl = nl_MultLoop_acc_50_nl[19:0];
  assign nl_MultLoop_acc_35_nl = conv_s2u_20_22(MultLoop_acc_50_nl) + ({(~ (data_rsci_idat[557:540]))
      , 4'b0000});
  assign MultLoop_acc_35_nl = nl_MultLoop_acc_35_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_26_nl = conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_152_nl)))
      + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_21_nl))) + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_2_nl)
      + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_14_nl)))
      + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_35_nl)));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_26_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_26_nl[17:0];
  assign nl_MultLoop_acc_54_nl = conv_s2s_20_21({(~ (data_rsci_idat[305:288])) ,
      2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[305:288]));
  assign MultLoop_acc_54_nl = nl_MultLoop_acc_54_nl[20:0];
  assign nl_MultLoop_acc_22_nl = conv_s2s_21_26(MultLoop_acc_54_nl) + ({(data_rsci_idat[305:288])
      , 8'b00000100});
  assign MultLoop_acc_22_nl = nl_MultLoop_acc_22_nl[25:0];
  assign nl_MultLoop_acc_153_nl = conv_s2s_12_13(data_rsci_idat[359:348]) + 13'b0000000000001;
  assign MultLoop_acc_153_nl = nl_MultLoop_acc_153_nl[12:0];
  assign nl_MultLoop_acc_56_nl = (~ (data_rsci_idat[359:342])) + conv_s2s_16_18({(MultLoop_acc_153_nl)
      , (data_rsci_idat[347:345])});
  assign MultLoop_acc_56_nl = nl_MultLoop_acc_56_nl[17:0];
  assign nl_MultLoop_acc_37_nl = conv_s2u_18_22(MultLoop_acc_56_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[359:342])) , 3'b001});
  assign MultLoop_acc_37_nl = nl_MultLoop_acc_37_nl[21:0];
  assign nl_MultLoop_acc_58_nl = conv_s2s_24_25({(~ (data_rsci_idat[377:360])) ,
      6'b000100}) + conv_s2s_20_25({(~ (data_rsci_idat[377:360])) , 2'b01}) + conv_s2s_18_25(~
      (data_rsci_idat[377:360]));
  assign MultLoop_acc_58_nl = nl_MultLoop_acc_58_nl[24:0];
  assign nl_MultLoop_acc_26_nl = conv_s2s_25_26(MultLoop_acc_58_nl) + ({(data_rsci_idat[377:360])
      , 8'b01000000});
  assign MultLoop_acc_26_nl = nl_MultLoop_acc_26_nl[25:0];
  assign nl_MultLoop_acc_154_nl =  -conv_s2s_10_11(data_rsci_idat[395:386]);
  assign MultLoop_acc_154_nl = nl_MultLoop_acc_154_nl[10:0];
  assign nl_MultLoop_acc_60_nl = ({(data_rsci_idat[395:378]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_154_nl)
      , (~ (data_rsci_idat[385:378]))});
  assign MultLoop_acc_60_nl = nl_MultLoop_acc_60_nl[19:0];
  assign nl_MultLoop_acc_61_nl = conv_s2s_23_24({(data_rsci_idat[395:378]) , 5'b00000})
      + conv_s2s_20_24(MultLoop_acc_60_nl);
  assign MultLoop_acc_61_nl = nl_MultLoop_acc_61_nl[23:0];
  assign nl_MultLoop_acc_155_nl = conv_s2u_16_18(readslicef_24_16_8((MultLoop_acc_61_nl)))
      + (~ (data_rsci_idat[395:378]));
  assign MultLoop_acc_155_nl = nl_MultLoop_acc_155_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_19_nl = conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_22_nl)))
      + conv_s2s_17_18(readslicef_22_17_5((MultLoop_acc_37_nl))) + conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_26_nl)))
      + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_155_nl)));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_19_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_19_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_nl = (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_25_nl)
      + (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_26_nl) + (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_19_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_nl[17:0];
  assign nl_res_rsci_d  = (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_30_nl)
      + (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_nl);

  function automatic [15:0] readslicef_18_16_2;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_18_16_2 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_18_17_1;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_18_17_1 = tmp[16:0];
  end
  endfunction


  function automatic [16:0] readslicef_19_17_2;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_19_17_2 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_19_18_1;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_19_18_1 = tmp[17:0];
  end
  endfunction


  function automatic [12:0] readslicef_20_13_7;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_20_13_7 = tmp[12:0];
  end
  endfunction


  function automatic [16:0] readslicef_20_17_3;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_20_17_3 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_20_18_2;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_20_18_2 = tmp[17:0];
  end
  endfunction


  function automatic [12:0] readslicef_21_13_8;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_21_13_8 = tmp[12:0];
  end
  endfunction


  function automatic [13:0] readslicef_21_14_7;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_21_14_7 = tmp[13:0];
  end
  endfunction


  function automatic [15:0] readslicef_21_16_5;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_21_16_5 = tmp[15:0];
  end
  endfunction


  function automatic [17:0] readslicef_21_18_3;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_21_18_3 = tmp[17:0];
  end
  endfunction


  function automatic [15:0] readslicef_22_16_6;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_22_16_6 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_22_17_5;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_22_17_5 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_22_18_4;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_22_18_4 = tmp[17:0];
  end
  endfunction


  function automatic [14:0] readslicef_23_15_8;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_23_15_8 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_23_16_7;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_23_16_7 = tmp[15:0];
  end
  endfunction


  function automatic [17:0] readslicef_23_18_5;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_23_18_5 = tmp[17:0];
  end
  endfunction


  function automatic [13:0] readslicef_24_14_10;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_24_14_10 = tmp[13:0];
  end
  endfunction


  function automatic [15:0] readslicef_24_16_8;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_24_16_8 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_24_17_7;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_24_17_7 = tmp[16:0];
  end
  endfunction


  function automatic [15:0] readslicef_25_16_9;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_25_16_9 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_25_17_8;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_25_17_8 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_25_18_7;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_25_18_7 = tmp[17:0];
  end
  endfunction


  function automatic [16:0] readslicef_26_17_9;
    input [25:0] vector;
    reg [25:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_26_17_9 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_26_18_8;
    input [25:0] vector;
    reg [25:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_26_18_8 = tmp[17:0];
  end
  endfunction


  function automatic [17:0] readslicef_28_18_10;
    input [27:0] vector;
    reg [27:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_28_18_10 = tmp[17:0];
  end
  endfunction


  function automatic [7:0] conv_s2s_7_8 ;
    input [6:0]  vector ;
  begin
    conv_s2s_7_8 = {vector[6], vector};
  end
  endfunction


  function automatic [8:0] conv_s2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_9 = {vector[7], vector};
  end
  endfunction


  function automatic [9:0] conv_s2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_10 = {vector[8], vector};
  end
  endfunction


  function automatic [10:0] conv_s2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_s2s_10_11 = {vector[9], vector};
  end
  endfunction


  function automatic [11:0] conv_s2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_12 = {vector[10], vector};
  end
  endfunction


  function automatic [12:0] conv_s2s_12_13 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_13 = {vector[11], vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_13_18 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_18 = {{5{vector[12]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_14_18 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_18 = {{4{vector[13]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_15_16 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_16 = {vector[14], vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_15_18 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_18 = {{3{vector[14]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_15_20 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_20 = {{5{vector[14]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_16_18 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_18 = {{2{vector[15]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_16_20 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_20 = {{4{vector[15]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_17_18 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_18 = {vector[16], vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_17_22 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_22 = {{5{vector[16]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_17_23 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_23 = {{6{vector[16]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_17_24 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_24 = {{7{vector[16]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_18_20 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_20 = {{2{vector[17]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_18_21 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_21 = {{3{vector[17]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_18_22 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_22 = {{4{vector[17]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_18_23 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_23 = {{5{vector[17]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_18_24 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_24 = {{6{vector[17]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_18_25 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_25 = {{7{vector[17]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_19_20 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_20 = {vector[18], vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_19_21 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_21 = {{2{vector[18]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_19_22 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_22 = {{3{vector[18]}}, vector};
  end
  endfunction


  function automatic [27:0] conv_s2s_19_28 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_28 = {{9{vector[18]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_20_21 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_21 = {vector[19], vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_20_22 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_22 = {{2{vector[19]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_20_23 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_23 = {{3{vector[19]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_20_24 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_24 = {{4{vector[19]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_20_25 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_25 = {{5{vector[19]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_21_23 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_23 = {{2{vector[20]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_21_24 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_24 = {{3{vector[20]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_21_26 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_26 = {{5{vector[20]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_22_23 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_23 = {vector[21], vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_22_24 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_24 = {{2{vector[21]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_22_25 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_25 = {{3{vector[21]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_23_24 ;
    input [22:0]  vector ;
  begin
    conv_s2s_23_24 = {vector[22], vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_24_25 ;
    input [23:0]  vector ;
  begin
    conv_s2s_24_25 = {vector[23], vector};
  end
  endfunction


  function automatic [27:0] conv_s2s_24_28 ;
    input [23:0]  vector ;
  begin
    conv_s2s_24_28 = {{4{vector[23]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_25_26 ;
    input [24:0]  vector ;
  begin
    conv_s2s_25_26 = {vector[24], vector};
  end
  endfunction


  function automatic [27:0] conv_s2s_27_28 ;
    input [26:0]  vector ;
  begin
    conv_s2s_27_28 = {vector[26], vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_13_18 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_18 = {{5{vector[12]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_14_18 ;
    input [13:0]  vector ;
  begin
    conv_s2u_14_18 = {{4{vector[13]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_14_19 ;
    input [13:0]  vector ;
  begin
    conv_s2u_14_19 = {{5{vector[13]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_15_18 ;
    input [14:0]  vector ;
  begin
    conv_s2u_15_18 = {{3{vector[14]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_15_19 ;
    input [14:0]  vector ;
  begin
    conv_s2u_15_19 = {{4{vector[14]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2u_16_17 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_17 = {vector[15], vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_16_18 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_18 = {{2{vector[15]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_16_19 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_19 = {{3{vector[15]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_17_18 ;
    input [16:0]  vector ;
  begin
    conv_s2u_17_18 = {vector[16], vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_17_19 ;
    input [16:0]  vector ;
  begin
    conv_s2u_17_19 = {{2{vector[16]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_19 = {vector[17], vector};
  end
  endfunction


  function automatic [19:0] conv_s2u_18_20 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_20 = {{2{vector[17]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2u_18_21 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_21 = {{3{vector[17]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_18_22 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_22 = {{4{vector[17]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2u_20_21 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_21 = {vector[19], vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_20_22 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_22 = {{2{vector[19]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_20_23 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_23 = {{3{vector[19]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_21_22 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_22 = {vector[20], vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_22_23 ;
    input [21:0]  vector ;
  begin
    conv_s2u_22_23 = {vector[21], vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_22_25 ;
    input [21:0]  vector ;
  begin
    conv_s2u_22_25 = {{3{vector[21]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_23_25 ;
    input [22:0]  vector ;
  begin
    conv_s2u_23_25 = {{2{vector[22]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2u_23_26 ;
    input [22:0]  vector ;
  begin
    conv_s2u_23_26 = {{3{vector[22]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_24_25 ;
    input [23:0]  vector ;
  begin
    conv_s2u_24_25 = {vector[23], vector};
  end
  endfunction


  function automatic [25:0] conv_s2u_25_26 ;
    input [24:0]  vector ;
  begin
    conv_s2u_25_26 = {vector[24], vector};
  end
  endfunction


  function automatic [15:0] conv_u2s_7_16 ;
    input [6:0]  vector ;
  begin
    conv_u2s_7_16 = {{9{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    nnet_dense_large_layer3_t_layer4_t_config4
// ------------------------------------------------------------------


module nnet_dense_large_layer3_t_layer4_t_config4 (
  data_rsc_dat, res_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_srst,
      ccs_ccore_en
);
  input [575:0] data_rsc_dat;
  output [17:0] res_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  nnet_dense_large_layer3_t_layer4_t_config4_core nnet_dense_large_layer3_t_layer4_t_config4_core_inst
      (
      .data_rsc_dat(data_rsc_dat),
      .res_rsc_z(res_rsc_z),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/nnet__relu_layer2_t_layer3_t_relu_config3__5caa6e7ac2e751923b640ab868b3dac817cc6_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4a/835166 Production Release
//  HLS Date:       Thu Sep  5 21:35:46 PDT 2019
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Mon Oct 21 13:59:59 2019
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    nnet_relu_layer2_t_layer3_t_relu_config3_core
// ------------------------------------------------------------------


module nnet_relu_layer2_t_layer3_t_relu_config3_core (
  data_rsc_dat, res_rsc_z, ccs_ccore_clk, ccs_ccore_srst, ccs_ccore_en
);
  input [575:0] data_rsc_dat;
  output [575:0] res_rsc_z;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [575:0] data_rsci_idat;
  reg [16:0] res_rsci_d_556_540;
  reg [16:0] res_rsci_d_538_522;
  reg [16:0] res_rsci_d_520_504;
  reg [16:0] res_rsci_d_502_486;
  reg [16:0] res_rsci_d_484_468;
  reg [16:0] res_rsci_d_466_450;
  reg [16:0] res_rsci_d_448_432;
  reg [16:0] res_rsci_d_430_414;
  reg [16:0] res_rsci_d_412_396;
  reg [16:0] res_rsci_d_394_378;
  reg [16:0] res_rsci_d_376_360;
  reg [16:0] res_rsci_d_358_342;
  reg [16:0] res_rsci_d_340_324;
  reg [16:0] res_rsci_d_322_306;
  reg [16:0] res_rsci_d_304_288;
  reg [16:0] res_rsci_d_286_270;
  reg [16:0] res_rsci_d_268_252;
  reg [16:0] res_rsci_d_250_234;
  reg [16:0] res_rsci_d_232_216;
  reg [16:0] res_rsci_d_214_198;
  reg [16:0] res_rsci_d_196_180;
  reg [16:0] res_rsci_d_178_162;
  reg [16:0] res_rsci_d_160_144;
  reg [16:0] res_rsci_d_142_126;
  reg [16:0] res_rsci_d_124_108;
  reg [16:0] res_rsci_d_106_90;
  reg [16:0] res_rsci_d_88_72;
  reg [16:0] res_rsci_d_70_54;
  reg [16:0] res_rsci_d_52_36;
  reg [16:0] res_rsci_d_34_18;
  reg [16:0] res_rsci_d_16_0;
  reg [16:0] res_rsci_d_574_558;

  wire[18:0] for_32_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_32_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_31_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_31_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_30_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_30_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_29_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_29_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_28_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_28_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_27_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_27_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_26_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_26_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_7_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_7_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_25_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_25_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_8_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_8_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_24_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_24_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_9_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_9_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_23_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_23_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_10_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_10_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_22_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_22_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_11_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_11_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_21_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_21_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_12_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_12_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_20_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_20_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_13_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_13_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_19_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_19_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_14_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_14_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_18_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_18_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_15_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_15_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_17_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_17_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_16_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_16_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [575:0] nl_res_rsci_d;
  assign nl_res_rsci_d = {1'b0 , res_rsci_d_574_558 , 1'b0 , res_rsci_d_556_540 ,
      1'b0 , res_rsci_d_538_522 , 1'b0 , res_rsci_d_520_504 , 1'b0 , res_rsci_d_502_486
      , 1'b0 , res_rsci_d_484_468 , 1'b0 , res_rsci_d_466_450 , 1'b0 , res_rsci_d_448_432
      , 1'b0 , res_rsci_d_430_414 , 1'b0 , res_rsci_d_412_396 , 1'b0 , res_rsci_d_394_378
      , 1'b0 , res_rsci_d_376_360 , 1'b0 , res_rsci_d_358_342 , 1'b0 , res_rsci_d_340_324
      , 1'b0 , res_rsci_d_322_306 , 1'b0 , res_rsci_d_304_288 , 1'b0 , res_rsci_d_286_270
      , 1'b0 , res_rsci_d_268_252 , 1'b0 , res_rsci_d_250_234 , 1'b0 , res_rsci_d_232_216
      , 1'b0 , res_rsci_d_214_198 , 1'b0 , res_rsci_d_196_180 , 1'b0 , res_rsci_d_178_162
      , 1'b0 , res_rsci_d_160_144 , 1'b0 , res_rsci_d_142_126 , 1'b0 , res_rsci_d_124_108
      , 1'b0 , res_rsci_d_106_90 , 1'b0 , res_rsci_d_88_72 , 1'b0 , res_rsci_d_70_54
      , 1'b0 , res_rsci_d_52_36 , 1'b0 , res_rsci_d_34_18 , 1'b0 , res_rsci_d_16_0};
  ccs_in_v1 #(.rscid(32'sd6),
  .width(32'sd576)) data_rsci (
      .dat(data_rsc_dat),
      .idat(data_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd7),
  .width(32'sd576)) res_rsci (
      .d(nl_res_rsci_d[575:0]),
      .z(res_rsc_z)
    );
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      res_rsci_d_574_558 <= 17'b00000000000000000;
      res_rsci_d_16_0 <= 17'b00000000000000000;
      res_rsci_d_556_540 <= 17'b00000000000000000;
      res_rsci_d_34_18 <= 17'b00000000000000000;
      res_rsci_d_538_522 <= 17'b00000000000000000;
      res_rsci_d_52_36 <= 17'b00000000000000000;
      res_rsci_d_520_504 <= 17'b00000000000000000;
      res_rsci_d_70_54 <= 17'b00000000000000000;
      res_rsci_d_502_486 <= 17'b00000000000000000;
      res_rsci_d_88_72 <= 17'b00000000000000000;
      res_rsci_d_484_468 <= 17'b00000000000000000;
      res_rsci_d_106_90 <= 17'b00000000000000000;
      res_rsci_d_466_450 <= 17'b00000000000000000;
      res_rsci_d_124_108 <= 17'b00000000000000000;
      res_rsci_d_448_432 <= 17'b00000000000000000;
      res_rsci_d_142_126 <= 17'b00000000000000000;
      res_rsci_d_430_414 <= 17'b00000000000000000;
      res_rsci_d_160_144 <= 17'b00000000000000000;
      res_rsci_d_412_396 <= 17'b00000000000000000;
      res_rsci_d_178_162 <= 17'b00000000000000000;
      res_rsci_d_394_378 <= 17'b00000000000000000;
      res_rsci_d_196_180 <= 17'b00000000000000000;
      res_rsci_d_376_360 <= 17'b00000000000000000;
      res_rsci_d_214_198 <= 17'b00000000000000000;
      res_rsci_d_358_342 <= 17'b00000000000000000;
      res_rsci_d_232_216 <= 17'b00000000000000000;
      res_rsci_d_340_324 <= 17'b00000000000000000;
      res_rsci_d_250_234 <= 17'b00000000000000000;
      res_rsci_d_322_306 <= 17'b00000000000000000;
      res_rsci_d_268_252 <= 17'b00000000000000000;
      res_rsci_d_304_288 <= 17'b00000000000000000;
      res_rsci_d_286_270 <= 17'b00000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      res_rsci_d_574_558 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[574:558]),
          (readslicef_19_1_18((for_32_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_16_0 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[16:0]),
          (readslicef_19_1_18((for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_556_540 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[556:540]),
          (readslicef_19_1_18((for_31_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_34_18 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[34:18]),
          (readslicef_19_1_18((for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_538_522 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[538:522]),
          (readslicef_19_1_18((for_30_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_52_36 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[52:36]),
          (readslicef_19_1_18((for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_520_504 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[520:504]),
          (readslicef_19_1_18((for_29_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_70_54 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[70:54]),
          (readslicef_19_1_18((for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_502_486 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[502:486]),
          (readslicef_19_1_18((for_28_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_88_72 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[88:72]),
          (readslicef_19_1_18((for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_484_468 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[484:468]),
          (readslicef_19_1_18((for_27_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_106_90 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[106:90]),
          (readslicef_19_1_18((for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_466_450 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[466:450]),
          (readslicef_19_1_18((for_26_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_124_108 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[124:108]),
          (readslicef_19_1_18((for_7_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_448_432 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[448:432]),
          (readslicef_19_1_18((for_25_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_142_126 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[142:126]),
          (readslicef_19_1_18((for_8_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_430_414 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[430:414]),
          (readslicef_19_1_18((for_24_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_160_144 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[160:144]),
          (readslicef_19_1_18((for_9_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_412_396 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[412:396]),
          (readslicef_19_1_18((for_23_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_178_162 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[178:162]),
          (readslicef_19_1_18((for_10_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_394_378 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[394:378]),
          (readslicef_19_1_18((for_22_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_196_180 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[196:180]),
          (readslicef_19_1_18((for_11_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_376_360 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[376:360]),
          (readslicef_19_1_18((for_21_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_214_198 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[214:198]),
          (readslicef_19_1_18((for_12_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_358_342 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[358:342]),
          (readslicef_19_1_18((for_20_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_232_216 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[232:216]),
          (readslicef_19_1_18((for_13_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_340_324 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[340:324]),
          (readslicef_19_1_18((for_19_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_250_234 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[250:234]),
          (readslicef_19_1_18((for_14_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_322_306 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[322:306]),
          (readslicef_19_1_18((for_18_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_268_252 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[268:252]),
          (readslicef_19_1_18((for_15_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_304_288 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[304:288]),
          (readslicef_19_1_18((for_17_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_286_270 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[286:270]),
          (readslicef_19_1_18((for_16_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
    end
  end
  assign nl_for_32_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[575:558]);
  assign for_32_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_32_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[17:0]);
  assign for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_31_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[557:540]);
  assign for_31_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_31_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[35:18]);
  assign for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_30_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[539:522]);
  assign for_30_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_30_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[53:36]);
  assign for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_29_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[521:504]);
  assign for_29_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_29_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[71:54]);
  assign for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_28_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[503:486]);
  assign for_28_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_28_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[89:72]);
  assign for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_27_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[485:468]);
  assign for_27_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_27_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[107:90]);
  assign for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_26_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[467:450]);
  assign for_26_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_26_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_7_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[125:108]);
  assign for_7_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_7_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_25_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[449:432]);
  assign for_25_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_25_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_8_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[143:126]);
  assign for_8_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_8_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_24_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[431:414]);
  assign for_24_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_24_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_9_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[161:144]);
  assign for_9_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_9_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_23_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[413:396]);
  assign for_23_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_23_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_10_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[179:162]);
  assign for_10_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_10_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_22_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[395:378]);
  assign for_22_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_22_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_11_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[197:180]);
  assign for_11_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_11_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_21_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[377:360]);
  assign for_21_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_21_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_12_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[215:198]);
  assign for_12_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_12_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_20_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[359:342]);
  assign for_20_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_20_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_13_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[233:216]);
  assign for_13_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_13_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_19_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[341:324]);
  assign for_19_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_19_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_14_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[251:234]);
  assign for_14_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_14_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_18_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[323:306]);
  assign for_18_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_18_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_15_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[269:252]);
  assign for_15_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_15_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_17_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[305:288]);
  assign for_17_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_17_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_16_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[287:270]);
  assign for_16_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_16_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];

  function automatic [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_19_1_18;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 18;
    readslicef_19_1_18 = tmp[0:0];
  end
  endfunction


  function automatic [18:0] conv_s2s_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_19 = {vector[17], vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    nnet_relu_layer2_t_layer3_t_relu_config3
// ------------------------------------------------------------------


module nnet_relu_layer2_t_layer3_t_relu_config3 (
  data_rsc_dat, res_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_srst,
      ccs_ccore_en
);
  input [575:0] data_rsc_dat;
  output [575:0] res_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  nnet_relu_layer2_t_layer3_t_relu_config3_core nnet_relu_layer2_t_layer3_t_relu_config3_core_inst
      (
      .data_rsc_dat(data_rsc_dat),
      .res_rsc_z(res_rsc_z),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/nnet__dense_large_input_t_layer2_t_config2__590166dd44e83a1ed2ecd69eb802a1da64c25_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4a/835166 Production Release
//  HLS Date:       Thu Sep  5 21:35:46 PDT 2019
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Mon Oct 21 14:02:23 2019
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    nnet_dense_large_input_t_layer2_t_config2_core
// ------------------------------------------------------------------


module nnet_dense_large_input_t_layer2_t_config2_core (
  data_rsc_dat, res_rsc_z, ccs_ccore_clk, ccs_ccore_srst, ccs_ccore_en
);
  input [179:0] data_rsc_dat;
  output [575:0] res_rsc_z;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [179:0] data_rsci_idat;
  reg [17:0] res_rsci_d_575_558;
  wire [18:0] nl_res_rsci_d_575_558;
  reg [17:0] res_rsci_d_557_540;
  wire [20:0] nl_res_rsci_d_557_540;
  reg [17:0] res_rsci_d_539_522;
  wire [20:0] nl_res_rsci_d_539_522;
  reg [17:0] res_rsci_d_521_504;
  wire [19:0] nl_res_rsci_d_521_504;
  reg [17:0] res_rsci_d_503_486;
  wire [18:0] nl_res_rsci_d_503_486;
  reg [17:0] res_rsci_d_485_468;
  wire [20:0] nl_res_rsci_d_485_468;
  reg [17:0] res_rsci_d_467_450;
  wire [20:0] nl_res_rsci_d_467_450;
  reg [17:0] res_rsci_d_449_432;
  wire [19:0] nl_res_rsci_d_449_432;
  reg [17:0] res_rsci_d_431_414;
  wire [20:0] nl_res_rsci_d_431_414;
  reg [17:0] res_rsci_d_413_396;
  wire [20:0] nl_res_rsci_d_413_396;
  reg [17:0] res_rsci_d_395_378;
  wire [19:0] nl_res_rsci_d_395_378;
  reg [17:0] res_rsci_d_377_360;
  wire [19:0] nl_res_rsci_d_377_360;
  reg [17:0] res_rsci_d_359_342;
  wire [20:0] nl_res_rsci_d_359_342;
  reg [17:0] res_rsci_d_341_324;
  wire [18:0] nl_res_rsci_d_341_324;
  reg [17:0] res_rsci_d_323_306;
  wire [18:0] nl_res_rsci_d_323_306;
  reg [17:0] res_rsci_d_305_288;
  wire [18:0] nl_res_rsci_d_305_288;
  reg [17:0] res_rsci_d_287_270;
  wire [20:0] nl_res_rsci_d_287_270;
  reg [17:0] res_rsci_d_269_252;
  wire [20:0] nl_res_rsci_d_269_252;
  reg [17:0] res_rsci_d_251_234;
  wire [20:0] nl_res_rsci_d_251_234;
  reg [17:0] res_rsci_d_233_216;
  wire [18:0] nl_res_rsci_d_233_216;
  reg [17:0] res_rsci_d_215_198;
  wire [18:0] nl_res_rsci_d_215_198;
  reg [17:0] res_rsci_d_197_180;
  wire [18:0] nl_res_rsci_d_197_180;
  reg [17:0] res_rsci_d_179_162;
  wire [18:0] nl_res_rsci_d_179_162;
  reg [17:0] res_rsci_d_161_144;
  wire [20:0] nl_res_rsci_d_161_144;
  reg [17:0] res_rsci_d_143_126;
  wire [19:0] nl_res_rsci_d_143_126;
  reg [17:0] res_rsci_d_125_108;
  wire [20:0] nl_res_rsci_d_125_108;
  reg [17:0] res_rsci_d_107_90;
  wire [18:0] nl_res_rsci_d_107_90;
  reg [17:0] res_rsci_d_89_72;
  wire [20:0] nl_res_rsci_d_89_72;
  reg [17:0] res_rsci_d_71_54;
  wire [18:0] nl_res_rsci_d_71_54;
  reg [17:0] res_rsci_d_53_36;
  wire [18:0] nl_res_rsci_d_53_36;
  reg [17:0] res_rsci_d_35_18;
  wire [18:0] nl_res_rsci_d_35_18;
  reg [17:0] res_rsci_d_17_0;
  wire [18:0] nl_res_rsci_d_17_0;
  wire [18:0] Result_acc_175_cse;
  wire [19:0] nl_Result_acc_175_cse;
  wire [20:0] MultLoop_acc_759_sdt_1;
  wire [21:0] nl_MultLoop_acc_759_sdt_1;
  wire [11:0] MultLoop_acc_1254_cse_1;
  wire [12:0] nl_MultLoop_acc_1254_cse_1;
  wire [8:0] MultLoop_acc_1213_cse_1;
  wire [9:0] nl_MultLoop_acc_1213_cse_1;
  wire [9:0] MultLoop_acc_1273_cse_1;
  wire [10:0] nl_MultLoop_acc_1273_cse_1;
  wire [18:0] MultLoop_acc_875_cse_1;
  wire [19:0] nl_MultLoop_acc_875_cse_1;
  wire [21:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_5_cse_1;
  wire [22:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_5_cse_1;
  wire [11:0] MultLoop_acc_1148_cse_1;
  wire [12:0] nl_MultLoop_acc_1148_cse_1;
  wire [17:0] MultLoop_acc_634_cse_1;
  wire [18:0] nl_MultLoop_acc_634_cse_1;
  wire [21:0] MultLoop_acc_839_cse_1;
  wire [22:0] nl_MultLoop_acc_839_cse_1;
  wire [19:0] MultLoop_acc_892_cse_1;
  wire [20:0] nl_MultLoop_acc_892_cse_1;
  wire [8:0] MultLoop_acc_1203_cse_1;
  wire [9:0] nl_MultLoop_acc_1203_cse_1;
  wire [20:0] MultLoop_acc_623_cse_1;
  wire [21:0] nl_MultLoop_acc_623_cse_1;
  wire [12:0] MultLoop_acc_1178_cse_1;
  wire [13:0] nl_MultLoop_acc_1178_cse_1;
  wire [20:0] MultLoop_acc_565_cse_1;
  wire [21:0] nl_MultLoop_acc_565_cse_1;
  wire [19:0] MultLoop_acc_777_sdt_1;
  wire [20:0] nl_MultLoop_acc_777_sdt_1;
  wire [11:0] Result_acc_207_cse_1;
  wire [12:0] nl_Result_acc_207_cse_1;
  wire [17:0] MultLoop_acc_543_cse_1;
  wire [18:0] nl_MultLoop_acc_543_cse_1;
  wire [17:0] MultLoop_acc_1017_cse_1;
  wire [18:0] nl_MultLoop_acc_1017_cse_1;
  wire [18:0] MultLoop_acc_405_cse_1;
  wire [19:0] nl_MultLoop_acc_405_cse_1;
  wire [21:0] MultLoop_acc_473_cse_1;
  wire [22:0] nl_MultLoop_acc_473_cse_1;
  wire [20:0] MultLoop_acc_763_cse_1;
  wire [21:0] nl_MultLoop_acc_763_cse_1;
  wire [9:0] Result_acc_202_cse_1;
  wire [10:0] nl_Result_acc_202_cse_1;
  wire [17:0] Result_acc_195_cse_1;
  wire [18:0] nl_Result_acc_195_cse_1;
  wire [18:0] MultLoop_acc_650_cse_1;
  wire [19:0] nl_MultLoop_acc_650_cse_1;
  wire [10:0] MultLoop_acc_1151_cse_1;
  wire [11:0] nl_MultLoop_acc_1151_cse_1;
  wire [17:0] MultLoop_acc_557_cse_1;
  wire [18:0] nl_MultLoop_acc_557_cse_1;
  wire [20:0] MultLoop_acc_789_cse_1;
  wire [21:0] nl_MultLoop_acc_789_cse_1;
  wire [17:0] MultLoop_acc_412_cse_1;
  wire [18:0] nl_MultLoop_acc_412_cse_1;
  wire [10:0] MultLoop_acc_1150_cse_1;
  wire [11:0] nl_MultLoop_acc_1150_cse_1;
  wire [17:0] MultLoop_acc_410_cse_1;
  wire [18:0] nl_MultLoop_acc_410_cse_1;
  wire [20:0] MultLoop_acc_744_cse_1;
  wire [21:0] nl_MultLoop_acc_744_cse_1;
  wire [19:0] MultLoop_acc_733_cse_1;
  wire [20:0] nl_MultLoop_acc_733_cse_1;
  wire [19:0] MultLoop_acc_805_cse_1;
  wire [20:0] nl_MultLoop_acc_805_cse_1;
  wire [18:0] MultLoop_acc_753_cse_1;
  wire [19:0] nl_MultLoop_acc_753_cse_1;
  wire [19:0] MultLoop_acc_786_cse_1;
  wire [20:0] nl_MultLoop_acc_786_cse_1;
  wire [20:0] MultLoop_acc_406_cse_1;
  wire [21:0] nl_MultLoop_acc_406_cse_1;
  wire [18:0] MultLoop_acc_812_cse_1;
  wire [19:0] nl_MultLoop_acc_812_cse_1;
  wire [17:0] MultLoop_acc_621_cse_1;
  wire [18:0] nl_MultLoop_acc_621_cse_1;
  wire [20:0] MultLoop_acc_399_cse_1;
  wire [21:0] nl_MultLoop_acc_399_cse_1;
  wire [21:0] MultLoop_acc_560_cse_1;
  wire [22:0] nl_MultLoop_acc_560_cse_1;
  wire [18:0] MultLoop_acc_702_cse_1;
  wire [19:0] nl_MultLoop_acc_702_cse_1;
  wire [20:0] MultLoop_acc_745_cse_1;
  wire [21:0] nl_MultLoop_acc_745_cse_1;
  wire [13:0] MultLoop_acc_1239_cse_1;
  wire [14:0] nl_MultLoop_acc_1239_cse_1;
  wire [17:0] MultLoop_acc_847_cse_1;
  wire [18:0] nl_MultLoop_acc_847_cse_1;
  wire [21:0] MultLoop_acc_578_cse_1;
  wire [22:0] nl_MultLoop_acc_578_cse_1;
  wire [17:0] MultLoop_acc_642_cse_1;
  wire [18:0] nl_MultLoop_acc_642_cse_1;
  wire [17:0] MultLoop_asn_361;
  wire [18:0] nl_MultLoop_asn_361;
  wire [9:0] Result_Result_conc_48_18_9;
  wire [10:0] nl_Result_Result_conc_48_18_9;
  wire [11:0] MultLoop_MultLoop_conc_202_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_202_18_7;
  wire [11:0] Result_Result_conc_50_13_2;
  wire [12:0] nl_Result_Result_conc_50_13_2;
  wire [9:0] MultLoop_MultLoop_conc_204_18_9;
  wire [10:0] nl_MultLoop_MultLoop_conc_204_18_9;
  wire [8:0] Result_Result_conc_52_18_10;
  wire [9:0] nl_Result_Result_conc_52_18_10;
  wire [10:0] Result_Result_conc_54_18_8;
  wire [11:0] nl_Result_Result_conc_54_18_8;
  wire [13:0] MultLoop_MultLoop_conc_206_18_5;
  wire [14:0] nl_MultLoop_MultLoop_conc_206_18_5;
  wire [10:0] MultLoop_MultLoop_conc_208_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_208_18_8;
  wire [12:0] Result_Result_conc_56_18_6;
  wire [13:0] nl_Result_Result_conc_56_18_6;
  wire [10:0] MultLoop_MultLoop_conc_210_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_210_18_8;
  wire [9:0] Result_Result_conc_58_18_9;
  wire [10:0] nl_Result_Result_conc_58_18_9;
  wire [12:0] MultLoop_MultLoop_conc_212_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_212_18_6;
  wire [8:0] MultLoop_MultLoop_conc_214_18_10;
  wire [9:0] nl_MultLoop_MultLoop_conc_214_18_10;
  wire [11:0] Result_Result_conc_60_18_7;
  wire [12:0] nl_Result_Result_conc_60_18_7;
  wire [10:0] MultLoop_MultLoop_conc_216_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_216_18_8;
  wire [12:0] Result_Result_conc_62_18_6;
  wire [13:0] nl_Result_Result_conc_62_18_6;
  wire [10:0] MultLoop_MultLoop_conc_218_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_218_18_8;
  wire [9:0] MultLoop_MultLoop_conc_222_18_9;
  wire [10:0] nl_MultLoop_MultLoop_conc_222_18_9;
  wire [10:0] MultLoop_MultLoop_conc_224_16_6;
  wire [11:0] nl_MultLoop_MultLoop_conc_224_16_6;
  wire [12:0] MultLoop_MultLoop_conc_226_16_4;
  wire [13:0] nl_MultLoop_MultLoop_conc_226_16_4;
  wire [9:0] MultLoop_MultLoop_conc_228_18_9;
  wire [10:0] nl_MultLoop_MultLoop_conc_228_18_9;
  wire [10:0] Result_Result_conc_64_18_8;
  wire [11:0] nl_Result_Result_conc_64_18_8;
  wire [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_4_itm_18_2_1;
  wire [16:0] MultLoop_acc_594_itm_18_2_1;
  wire [10:0] Result_acc_71_itm_17_7;
  wire [16:0] MultLoop_acc_19_itm_19_3;
  wire [15:0] MultLoop_acc_213_itm_22_7;
  wire [13:0] Result_acc_46_itm_17_4;
  wire [15:0] MultLoop_acc_123_itm_21_6;
  wire [12:0] Result_acc_41_itm_20_8;
  wire [16:0] MultLoop_acc_302_itm_23_7;
  wire [13:0] MultLoop_acc_45_itm_22_9;
  wire [18:0] MultLoop_acc_808_itm_20_2_1;
  wire [16:0] MultLoop_acc_56_itm_17_1;
  wire [16:0] MultLoop_acc_74_itm_17_1;
  wire [15:0] MultLoop_acc_596_itm_20_5;
  wire [15:0] MultLoop_acc_714_itm_19_4;
  wire [14:0] MultLoop_acc_279_itm_20_6;
  wire [15:0] MultLoop_acc_916_itm_18_3;
  wire [17:0] MultLoop_acc_694_itm_19_2_1;
  wire [17:0] MultLoop_acc_1374_itm_18_1;
  wire [13:0] MultLoop_acc_237_itm_22_9;
  wire [16:0] MultLoop_acc_1354_itm_19_3;
  wire [16:0] MultLoop_acc_114_itm_19_3;
  wire [13:0] MultLoop_acc_108_itm_19_6;
  wire [16:0] MultLoop_acc_100_itm_23_7;
  wire [18:0] MultLoop_acc_554_itm_23_5_1;
  wire [17:0] MultLoop_acc_901_itm_22_5;
  wire [16:0] MultLoop_acc_751_itm_18_2;
  wire [15:0] MultLoop_acc_620_itm_18_3;
  wire [10:0] MultLoop_acc_130_itm_20_10;
  wire [14:0] MultLoop_acc_731_itm_18_4;
  wire [18:0] MultLoop_acc_660_itm_22_4_1;
  wire [16:0] MultLoop_acc_206_itm_20_4;
  wire [16:0] MultLoop_acc_1198_itm_18_2;
  wire [15:0] MultLoop_acc_159_itm_24_9;
  wire [9:0] MultLoop_acc_170_itm_17_8;
  wire [17:0] MultLoop_acc_1395_itm_20_3_1;
  wire [18:0] MultLoop_acc_1397_itm_21_3_1;
  wire [15:0] MultLoop_acc_1399_itm_20_5;
  wire [15:0] MultLoop_acc_1401_itm_20_5;
  wire [18:0] MultLoop_acc_1403_itm_20_2_1;
  wire [15:0] MultLoop_acc_1348_itm_18_3;
  wire [13:0] MultLoop_acc_1350_itm_18_5;
  wire [16:0] MultLoop_acc_353_itm_22_6;
  wire [18:0] MultLoop_acc_1390_itm_22_4_1;
  wire [18:0] MultLoop_acc_1359_itm_20_2_1;

  wire[17:0] MultLoop_acc_421_nl;
  wire[18:0] nl_MultLoop_acc_421_nl;
  wire[17:0] MultLoop_acc_419_nl;
  wire[18:0] nl_MultLoop_acc_419_nl;
  wire[20:0] Result_acc_242_nl;
  wire[21:0] nl_Result_acc_242_nl;
  wire[25:0] Result_acc_94_nl;
  wire[26:0] nl_Result_acc_94_nl;
  wire[16:0] MultLoop_acc_416_nl;
  wire[17:0] nl_MultLoop_acc_416_nl;
  wire[24:0] Result_acc_70_nl;
  wire[25:0] nl_Result_acc_70_nl;
  wire[22:0] Result_acc_87_nl;
  wire[23:0] nl_Result_acc_87_nl;
  wire[17:0] Result_acc_244_nl;
  wire[18:0] nl_Result_acc_244_nl;
  wire[23:0] Result_acc_90_nl;
  wire[25:0] nl_Result_acc_90_nl;
  wire[16:0] MultLoop_acc_418_nl;
  wire[17:0] nl_MultLoop_acc_418_nl;
  wire[15:0] MultLoop_acc_415_nl;
  wire[16:0] nl_MultLoop_acc_415_nl;
  wire[13:0] MultLoop_acc_414_nl;
  wire[14:0] nl_MultLoop_acc_414_nl;
  wire[8:0] MultLoop_acc_1347_nl;
  wire[9:0] nl_MultLoop_acc_1347_nl;
  wire[17:0] MultLoop_acc_420_nl;
  wire[18:0] nl_MultLoop_acc_420_nl;
  wire[17:0] MultLoop_acc_417_nl;
  wire[18:0] nl_MultLoop_acc_417_nl;
  wire[17:0] Result_acc_246_nl;
  wire[18:0] nl_Result_acc_246_nl;
  wire[21:0] Result_acc_92_nl;
  wire[22:0] nl_Result_acc_92_nl;
  wire[21:0] Result_acc_79_nl;
  wire[22:0] nl_Result_acc_79_nl;
  wire[17:0] Result_acc_85_nl;
  wire[18:0] nl_Result_acc_85_nl;
  wire[17:0] MultLoop_acc_1146_nl;
  wire[18:0] nl_MultLoop_acc_1146_nl;
  wire[17:0] MultLoop_acc_1144_nl;
  wire[18:0] nl_MultLoop_acc_1144_nl;
  wire[22:0] MultLoop_acc_16_nl;
  wire[23:0] nl_MultLoop_acc_16_nl;
  wire[18:0] MultLoop_acc_1136_nl;
  wire[19:0] nl_MultLoop_acc_1136_nl;
  wire[18:0] MultLoop_acc_294_nl;
  wire[19:0] nl_MultLoop_acc_294_nl;
  wire[17:0] MultLoop_acc_1143_nl;
  wire[20:0] nl_MultLoop_acc_1143_nl;
  wire[21:0] MultLoop_acc_12_nl;
  wire[22:0] nl_MultLoop_acc_12_nl;
  wire[13:0] MultLoop_acc_1138_nl;
  wire[14:0] nl_MultLoop_acc_1138_nl;
  wire[19:0] MultLoop_acc_18_nl;
  wire[20:0] nl_MultLoop_acc_18_nl;
  wire[9:0] MultLoop_acc_1343_nl;
  wire[10:0] nl_MultLoop_acc_1343_nl;
  wire[19:0] MultLoop_acc_293_nl;
  wire[20:0] nl_MultLoop_acc_293_nl;
  wire[17:0] MultLoop_acc_1124_nl;
  wire[18:0] nl_MultLoop_acc_1124_nl;
  wire[17:0] MultLoop_acc_1145_nl;
  wire[18:0] nl_MultLoop_acc_1145_nl;
  wire[17:0] MultLoop_acc_1142_nl;
  wire[18:0] nl_MultLoop_acc_1142_nl;
  wire[22:0] MultLoop_acc_22_nl;
  wire[23:0] nl_MultLoop_acc_22_nl;
  wire[20:0] MultLoop_acc_1127_nl;
  wire[22:0] nl_MultLoop_acc_1127_nl;
  wire[24:0] MultLoop_acc_292_nl;
  wire[25:0] nl_MultLoop_acc_292_nl;
  wire[19:0] MultLoop_acc_1129_nl;
  wire[20:0] nl_MultLoop_acc_1129_nl;
  wire[19:0] MultLoop_acc_1346_nl;
  wire[20:0] nl_MultLoop_acc_1346_nl;
  wire[26:0] MultLoop_acc_1134_nl;
  wire[28:0] nl_MultLoop_acc_1134_nl;
  wire[21:0] MultLoop_acc_1132_nl;
  wire[22:0] nl_MultLoop_acc_1132_nl;
  wire[19:0] MultLoop_acc_1131_nl;
  wire[20:0] nl_MultLoop_acc_1131_nl;
  wire[17:0] MultLoop_acc_429_nl;
  wire[19:0] nl_MultLoop_acc_429_nl;
  wire[17:0] Result_acc_237_nl;
  wire[18:0] nl_Result_acc_237_nl;
  wire[22:0] Result_acc_108_nl;
  wire[23:0] nl_Result_acc_108_nl;
  wire[19:0] Result_acc_107_nl;
  wire[20:0] nl_Result_acc_107_nl;
  wire[17:0] Result_acc_106_nl;
  wire[18:0] nl_Result_acc_106_nl;
  wire[9:0] Result_acc_236_nl;
  wire[10:0] nl_Result_acc_236_nl;
  wire[26:0] Result_acc_60_nl;
  wire[27:0] nl_Result_acc_60_nl;
  wire[17:0] Result_acc_239_nl;
  wire[18:0] nl_Result_acc_239_nl;
  wire[19:0] Result_acc_110_nl;
  wire[20:0] nl_Result_acc_110_nl;
  wire[25:0] Result_acc_63_nl;
  wire[27:0] nl_Result_acc_63_nl;
  wire[11:0] Result_acc_240_nl;
  wire[12:0] nl_Result_acc_240_nl;
  wire[17:0] MultLoop_acc_428_nl;
  wire[18:0] nl_MultLoop_acc_428_nl;
  wire[17:0] MultLoop_acc_424_nl;
  wire[18:0] nl_MultLoop_acc_424_nl;
  wire[26:0] Result_acc_64_nl;
  wire[27:0] nl_Result_acc_64_nl;
  wire[23:0] Result_acc_115_nl;
  wire[25:0] nl_Result_acc_115_nl;
  wire[20:0] Result_acc_66_nl;
  wire[21:0] nl_Result_acc_66_nl;
  wire[17:0] Result_acc_96_nl;
  wire[18:0] nl_Result_acc_96_nl;
  wire[18:0] Result_acc_232_nl;
  wire[19:0] nl_Result_acc_232_nl;
  wire[19:0] Result_acc_248_nl;
  wire[20:0] nl_Result_acc_248_nl;
  wire[16:0] MultLoop_acc_422_nl;
  wire[17:0] nl_MultLoop_acc_422_nl;
  wire[22:0] Result_acc_68_nl;
  wire[23:0] nl_Result_acc_68_nl;
  wire[20:0] Result_acc_104_nl;
  wire[21:0] nl_Result_acc_104_nl;
  wire[20:0] Result_acc_67_nl;
  wire[21:0] nl_Result_acc_67_nl;
  wire[17:0] Result_acc_98_nl;
  wire[18:0] nl_Result_acc_98_nl;
  wire[21:0] Result_acc_62_nl;
  wire[22:0] nl_Result_acc_62_nl;
  wire[20:0] Result_acc_101_nl;
  wire[22:0] nl_Result_acc_101_nl;
  wire[12:0] Result_acc_234_nl;
  wire[13:0] nl_Result_acc_234_nl;
  wire[17:0] MultLoop_acc_1123_nl;
  wire[18:0] nl_MultLoop_acc_1123_nl;
  wire[17:0] MultLoop_acc_1121_nl;
  wire[19:0] nl_MultLoop_acc_1121_nl;
  wire[18:0] MultLoop_acc_1330_nl;
  wire[19:0] nl_MultLoop_acc_1330_nl;
  wire[20:0] MultLoop_acc_296_nl;
  wire[21:0] nl_MultLoop_acc_296_nl;
  wire[18:0] MultLoop_acc_1098_nl;
  wire[19:0] nl_MultLoop_acc_1098_nl;
  wire[17:0] MultLoop_acc_1332_nl;
  wire[18:0] nl_MultLoop_acc_1332_nl;
  wire[24:0] MultLoop_acc_1101_nl;
  wire[25:0] nl_MultLoop_acc_1101_nl;
  wire[21:0] MultLoop_acc_1100_nl;
  wire[22:0] nl_MultLoop_acc_1100_nl;
  wire[10:0] MultLoop_acc_1331_nl;
  wire[11:0] nl_MultLoop_acc_1331_nl;
  wire[15:0] MultLoop_acc_1115_nl;
  wire[16:0] nl_MultLoop_acc_1115_nl;
  wire[17:0] MultLoop_acc_1334_nl;
  wire[18:0] nl_MultLoop_acc_1334_nl;
  wire[23:0] MultLoop_acc_1093_nl;
  wire[24:0] nl_MultLoop_acc_1093_nl;
  wire[10:0] MultLoop_acc_1333_nl;
  wire[11:0] nl_MultLoop_acc_1333_nl;
  wire[17:0] MultLoop_acc_1120_nl;
  wire[18:0] nl_MultLoop_acc_1120_nl;
  wire[27:0] MultLoop_acc_24_nl;
  wire[28:0] nl_MultLoop_acc_24_nl;
  wire[24:0] MultLoop_acc_1103_nl;
  wire[25:0] nl_MultLoop_acc_1103_nl;
  wire[17:0] MultLoop_acc_1337_nl;
  wire[18:0] nl_MultLoop_acc_1337_nl;
  wire[18:0] MultLoop_acc_1336_nl;
  wire[19:0] nl_MultLoop_acc_1336_nl;
  wire[22:0] MultLoop_acc_1106_nl;
  wire[24:0] nl_MultLoop_acc_1106_nl;
  wire[17:0] MultLoop_acc_1122_nl;
  wire[18:0] nl_MultLoop_acc_1122_nl;
  wire[17:0] MultLoop_acc_1119_nl;
  wire[18:0] nl_MultLoop_acc_1119_nl;
  wire[17:0] MultLoop_acc_1339_nl;
  wire[18:0] nl_MultLoop_acc_1339_nl;
  wire[22:0] MultLoop_acc_1110_nl;
  wire[24:0] nl_MultLoop_acc_1110_nl;
  wire[10:0] MultLoop_acc_1338_nl;
  wire[11:0] nl_MultLoop_acc_1338_nl;
  wire[23:0] MultLoop_acc_29_nl;
  wire[24:0] nl_MultLoop_acc_29_nl;
  wire[20:0] MultLoop_acc_1111_nl;
  wire[21:0] nl_MultLoop_acc_1111_nl;
  wire[17:0] MultLoop_acc_1118_nl;
  wire[18:0] nl_MultLoop_acc_1118_nl;
  wire[25:0] MultLoop_acc_297_nl;
  wire[26:0] nl_MultLoop_acc_297_nl;
  wire[20:0] MultLoop_acc_1114_nl;
  wire[21:0] nl_MultLoop_acc_1114_nl;
  wire[17:0] MultLoop_acc_1113_nl;
  wire[18:0] nl_MultLoop_acc_1113_nl;
  wire[19:0] MultLoop_acc_1341_nl;
  wire[20:0] nl_MultLoop_acc_1341_nl;
  wire[25:0] MultLoop_acc_1096_nl;
  wire[26:0] nl_MultLoop_acc_1096_nl;
  wire[22:0] MultLoop_acc_1095_nl;
  wire[23:0] nl_MultLoop_acc_1095_nl;
  wire[17:0] MultLoop_acc_439_nl;
  wire[18:0] nl_MultLoop_acc_439_nl;
  wire[17:0] MultLoop_acc_437_nl;
  wire[18:0] nl_MultLoop_acc_437_nl;
  wire[16:0] MultLoop_acc_433_nl;
  wire[17:0] nl_MultLoop_acc_433_nl;
  wire[21:0] Result_acc_55_nl;
  wire[22:0] nl_Result_acc_55_nl;
  wire[17:0] Result_acc_128_nl;
  wire[18:0] nl_Result_acc_128_nl;
  wire[12:0] Result_acc_223_nl;
  wire[13:0] nl_Result_acc_223_nl;
  wire[18:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_15_nl;
  wire[19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_15_nl;
  wire[20:0] Result_acc_226_nl;
  wire[21:0] nl_Result_acc_226_nl;
  wire[17:0] Result_acc_225_nl;
  wire[18:0] nl_Result_acc_225_nl;
  wire[22:0] Result_acc_130_nl;
  wire[23:0] nl_Result_acc_130_nl;
  wire[9:0] Result_acc_224_nl;
  wire[10:0] nl_Result_acc_224_nl;
  wire[17:0] MultLoop_acc_436_nl;
  wire[18:0] nl_MultLoop_acc_436_nl;
  wire[26:0] Result_acc_47_nl;
  wire[28:0] nl_Result_acc_47_nl;
  wire[21:0] Result_acc_251_nl;
  wire[22:0] nl_Result_acc_251_nl;
  wire[23:0] Result_acc_54_nl;
  wire[24:0] nl_Result_acc_54_nl;
  wire[22:0] Result_acc_121_nl;
  wire[23:0] nl_Result_acc_121_nl;
  wire[19:0] Result_acc_120_nl;
  wire[21:0] nl_Result_acc_120_nl;
  wire[22:0] Result_acc_53_nl;
  wire[23:0] nl_Result_acc_53_nl;
  wire[20:0] Result_acc_118_nl;
  wire[21:0] nl_Result_acc_118_nl;
  wire[12:0] MultLoop_acc_1329_nl;
  wire[13:0] nl_MultLoop_acc_1329_nl;
  wire[25:0] Result_acc_49_nl;
  wire[27:0] nl_Result_acc_49_nl;
  wire[17:0] Result_acc_230_nl;
  wire[18:0] nl_Result_acc_230_nl;
  wire[21:0] Result_acc_126_nl;
  wire[22:0] nl_Result_acc_126_nl;
  wire[10:0] Result_acc_229_nl;
  wire[11:0] nl_Result_acc_229_nl;
  wire[17:0] MultLoop_acc_1091_nl;
  wire[20:0] nl_MultLoop_acc_1091_nl;
  wire[17:0] MultLoop_acc_1324_nl;
  wire[18:0] nl_MultLoop_acc_1324_nl;
  wire[24:0] MultLoop_acc_1078_nl;
  wire[26:0] nl_MultLoop_acc_1078_nl;
  wire[14:0] MultLoop_acc_1085_nl;
  wire[15:0] nl_MultLoop_acc_1085_nl;
  wire[18:0] MultLoop_acc_1385_nl;
  wire[19:0] nl_MultLoop_acc_1385_nl;
  wire[23:0] MultLoop_acc_44_nl;
  wire[25:0] nl_MultLoop_acc_44_nl;
  wire[13:0] MultLoop_acc_1325_nl;
  wire[14:0] nl_MultLoop_acc_1325_nl;
  wire[14:0] MultLoop_22_MultLoop_acc_3_nl;
  wire[15:0] nl_MultLoop_22_MultLoop_acc_3_nl;
  wire[10:0] MultLoop_acc_34_nl;
  wire[11:0] nl_MultLoop_acc_34_nl;
  wire[20:0] MultLoop_acc_298_nl;
  wire[21:0] nl_MultLoop_acc_298_nl;
  wire[17:0] MultLoop_acc_1069_nl;
  wire[18:0] nl_MultLoop_acc_1069_nl;
  wire[13:0] MultLoop_acc_1326_nl;
  wire[14:0] nl_MultLoop_acc_1326_nl;
  wire[20:0] MultLoop_acc_299_nl;
  wire[21:0] nl_MultLoop_acc_299_nl;
  wire[18:0] MultLoop_acc_1072_nl;
  wire[19:0] nl_MultLoop_acc_1072_nl;
  wire[17:0] MultLoop_acc_1322_nl;
  wire[18:0] nl_MultLoop_acc_1322_nl;
  wire[22:0] MultLoop_acc_1074_nl;
  wire[23:0] nl_MultLoop_acc_1074_nl;
  wire[17:0] MultLoop_acc_1090_nl;
  wire[18:0] nl_MultLoop_acc_1090_nl;
  wire[25:0] MultLoop_acc_37_nl;
  wire[26:0] nl_MultLoop_acc_37_nl;
  wire[23:0] MultLoop_acc_1081_nl;
  wire[24:0] nl_MultLoop_acc_1081_nl;
  wire[17:0] MultLoop_acc_1080_nl;
  wire[18:0] nl_MultLoop_acc_1080_nl;
  wire[19:0] MultLoop_acc_1328_nl;
  wire[20:0] nl_MultLoop_acc_1328_nl;
  wire[26:0] MultLoop_acc_1084_nl;
  wire[27:0] nl_MultLoop_acc_1084_nl;
  wire[22:0] MultLoop_acc_1083_nl;
  wire[23:0] nl_MultLoop_acc_1083_nl;
  wire[17:0] MultLoop_acc_447_nl;
  wire[18:0] nl_MultLoop_acc_447_nl;
  wire[17:0] MultLoop_acc_444_nl;
  wire[18:0] nl_MultLoop_acc_444_nl;
  wire[24:0] Result_acc_37_nl;
  wire[26:0] nl_Result_acc_37_nl;
  wire[23:0] Result_acc_40_nl;
  wire[24:0] nl_Result_acc_40_nl;
  wire[22:0] Result_acc_146_nl;
  wire[23:0] nl_Result_acc_146_nl;
  wire[19:0] Result_acc_44_nl;
  wire[20:0] nl_Result_acc_44_nl;
  wire[17:0] Result_acc_147_nl;
  wire[18:0] nl_Result_acc_147_nl;
  wire[17:0] MultLoop_acc_446_nl;
  wire[18:0] nl_MultLoop_acc_446_nl;
  wire[18:0] Result_acc_217_nl;
  wire[19:0] nl_Result_acc_217_nl;
  wire[23:0] Result_acc_148_nl;
  wire[24:0] nl_Result_acc_148_nl;
  wire[16:0] MultLoop_acc_443_nl;
  wire[17:0] nl_MultLoop_acc_443_nl;
  wire[14:0] MultLoop_acc_442_nl;
  wire[16:0] nl_MultLoop_acc_442_nl;
  wire[11:0] MultLoop_acc_1320_nl;
  wire[12:0] nl_MultLoop_acc_1320_nl;
  wire[17:0] Result_acc_35_nl;
  wire[18:0] nl_Result_acc_35_nl;
  wire[18:0] Result_acc_42_nl;
  wire[19:0] nl_Result_acc_42_nl;
  wire[20:0] Result_acc_43_nl;
  wire[21:0] nl_Result_acc_43_nl;
  wire[17:0] Result_acc_140_nl;
  wire[18:0] nl_Result_acc_140_nl;
  wire[26:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_nl;
  wire[27:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_nl;
  wire[23:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_6_nl;
  wire[24:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_6_nl;
  wire[17:0] Result_acc_221_nl;
  wire[18:0] nl_Result_acc_221_nl;
  wire[19:0] Result_acc_142_nl;
  wire[20:0] nl_Result_acc_142_nl;
  wire[11:0] Result_acc_220_nl;
  wire[12:0] nl_Result_acc_220_nl;
  wire[17:0] MultLoop_acc_1065_nl;
  wire[19:0] nl_MultLoop_acc_1065_nl;
  wire[17:0] MultLoop_acc_1063_nl;
  wire[19:0] nl_MultLoop_acc_1063_nl;
  wire[22:0] MultLoop_acc_305_nl;
  wire[23:0] nl_MultLoop_acc_305_nl;
  wire[20:0] MultLoop_acc_1045_nl;
  wire[21:0] nl_MultLoop_acc_1045_nl;
  wire[17:0] MultLoop_acc_1044_nl;
  wire[18:0] nl_MultLoop_acc_1044_nl;
  wire[22:0] MultLoop_acc_53_nl;
  wire[23:0] nl_MultLoop_acc_53_nl;
  wire[20:0] MultLoop_acc_1047_nl;
  wire[21:0] nl_MultLoop_acc_1047_nl;
  wire[13:0] MultLoop_acc_1317_nl;
  wire[14:0] nl_MultLoop_acc_1317_nl;
  wire[16:0] MultLoop_34_MultLoop_acc_3_nl;
  wire[18:0] nl_MultLoop_34_MultLoop_acc_3_nl;
  wire[19:0] MultLoop_acc_1412_nl;
  wire[20:0] nl_MultLoop_acc_1412_nl;
  wire[10:0] MultLoop_acc_1319_nl;
  wire[11:0] nl_MultLoop_acc_1319_nl;
  wire[20:0] MultLoop_acc_1405_nl;
  wire[21:0] nl_MultLoop_acc_1405_nl;
  wire[19:0] MultLoop_acc_306_nl;
  wire[20:0] nl_MultLoop_acc_306_nl;
  wire[17:0] MultLoop_acc_1042_nl;
  wire[18:0] nl_MultLoop_acc_1042_nl;
  wire[17:0] MultLoop_acc_1064_nl;
  wire[18:0] nl_MultLoop_acc_1064_nl;
  wire[23:0] MultLoop_acc_303_nl;
  wire[24:0] nl_MultLoop_acc_303_nl;
  wire[22:0] MultLoop_acc_1058_nl;
  wire[24:0] nl_MultLoop_acc_1058_nl;
  wire[23:0] MultLoop_acc_304_nl;
  wire[24:0] nl_MultLoop_acc_304_nl;
  wire[21:0] MultLoop_acc_1060_nl;
  wire[22:0] nl_MultLoop_acc_1060_nl;
  wire[17:0] MultLoop_acc_457_nl;
  wire[18:0] nl_MultLoop_acc_457_nl;
  wire[17:0] MultLoop_acc_455_nl;
  wire[18:0] nl_MultLoop_acc_455_nl;
  wire[24:0] Result_acc_23_nl;
  wire[25:0] nl_Result_acc_23_nl;
  wire[23:0] Result_acc_162_nl;
  wire[24:0] nl_Result_acc_162_nl;
  wire[26:0] Result_acc_28_nl;
  wire[28:0] nl_Result_acc_28_nl;
  wire[17:0] MultLoop_acc_454_nl;
  wire[19:0] nl_MultLoop_acc_454_nl;
  wire[19:0] Result_acc_213_nl;
  wire[20:0] nl_Result_acc_213_nl;
  wire[17:0] Result_acc_212_nl;
  wire[18:0] nl_Result_acc_212_nl;
  wire[21:0] Result_acc_155_nl;
  wire[22:0] nl_Result_acc_155_nl;
  wire[17:0] Result_acc_25_nl;
  wire[18:0] nl_Result_acc_25_nl;
  wire[24:0] Result_acc_24_nl;
  wire[26:0] nl_Result_acc_24_nl;
  wire[17:0] MultLoop_acc_456_nl;
  wire[18:0] nl_MultLoop_acc_456_nl;
  wire[17:0] MultLoop_acc_453_nl;
  wire[19:0] nl_MultLoop_acc_453_nl;
  wire[21:0] Result_acc_27_nl;
  wire[22:0] nl_Result_acc_27_nl;
  wire[18:0] Result_acc_158_nl;
  wire[19:0] nl_Result_acc_158_nl;
  wire[22:0] Result_acc_31_nl;
  wire[23:0] nl_Result_acc_31_nl;
  wire[21:0] Result_acc_154_nl;
  wire[22:0] nl_Result_acc_154_nl;
  wire[11:0] MultLoop_acc_450_nl;
  wire[12:0] nl_MultLoop_acc_450_nl;
  wire[10:0] MultLoop_acc_449_nl;
  wire[11:0] nl_MultLoop_acc_449_nl;
  wire[20:0] Result_acc_21_nl;
  wire[21:0] nl_Result_acc_21_nl;
  wire[16:0] Result_acc_215_nl;
  wire[17:0] nl_Result_acc_215_nl;
  wire[24:0] Result_acc_32_nl;
  wire[25:0] nl_Result_acc_32_nl;
  wire[17:0] Result_acc_160_nl;
  wire[18:0] nl_Result_acc_160_nl;
  wire[17:0] MultLoop_acc_1040_nl;
  wire[19:0] nl_MultLoop_acc_1040_nl;
  wire[18:0] MultLoop_acc_1313_nl;
  wire[19:0] nl_MultLoop_acc_1313_nl;
  wire[21:0] MultLoop_acc_1384_nl;
  wire[22:0] nl_MultLoop_acc_1384_nl;
  wire[17:0] MultLoop_acc_1315_nl;
  wire[18:0] nl_MultLoop_acc_1315_nl;
  wire[23:0] MultLoop_acc_1030_nl;
  wire[25:0] nl_MultLoop_acc_1030_nl;
  wire[15:0] MultLoop_acc_57_nl;
  wire[16:0] nl_MultLoop_acc_57_nl;
  wire[20:0] MultLoop_acc_310_nl;
  wire[21:0] nl_MultLoop_acc_310_nl;
  wire[17:0] MultLoop_acc_1016_nl;
  wire[18:0] nl_MultLoop_acc_1016_nl;
  wire[17:0] MultLoop_acc_1039_nl;
  wire[18:0] nl_MultLoop_acc_1039_nl;
  wire[23:0] MultLoop_acc_309_nl;
  wire[24:0] nl_MultLoop_acc_309_nl;
  wire[21:0] MultLoop_acc_1033_nl;
  wire[22:0] nl_MultLoop_acc_1033_nl;
  wire[17:0] MultLoop_acc_1032_nl;
  wire[18:0] nl_MultLoop_acc_1032_nl;
  wire[11:0] MultLoop_acc_1309_nl;
  wire[12:0] nl_MultLoop_acc_1309_nl;
  wire[16:0] MultLoop_acc_1035_nl;
  wire[17:0] nl_MultLoop_acc_1035_nl;
  wire[20:0] MultLoop_acc_308_nl;
  wire[21:0] nl_MultLoop_acc_308_nl;
  wire[19:0] MultLoop_acc_60_nl;
  wire[20:0] nl_MultLoop_acc_60_nl;
  wire[18:0] MultLoop_acc_1019_nl;
  wire[19:0] nl_MultLoop_acc_1019_nl;
  wire[14:0] MultLoop_acc_1310_nl;
  wire[15:0] nl_MultLoop_acc_1310_nl;
  wire[18:0] MultLoop_acc_1312_nl;
  wire[19:0] nl_MultLoop_acc_1312_nl;
  wire[23:0] MultLoop_acc_1024_nl;
  wire[24:0] nl_MultLoop_acc_1024_nl;
  wire[21:0] MultLoop_acc_1023_nl;
  wire[22:0] nl_MultLoop_acc_1023_nl;
  wire[21:0] MultLoop_acc_307_nl;
  wire[22:0] nl_MultLoop_acc_307_nl;
  wire[20:0] MultLoop_acc_1021_nl;
  wire[21:0] nl_MultLoop_acc_1021_nl;
  wire[24:0] MultLoop_acc_65_nl;
  wire[26:0] nl_MultLoop_acc_65_nl;
  wire[17:0] MultLoop_acc_465_nl;
  wire[18:0] nl_MultLoop_acc_465_nl;
  wire[17:0] MultLoop_acc_462_nl;
  wire[18:0] nl_MultLoop_acc_462_nl;
  wire[20:0] Result_acc_252_nl;
  wire[21:0] nl_Result_acc_252_nl;
  wire[21:0] Result_acc_9_nl;
  wire[22:0] nl_Result_acc_9_nl;
  wire[18:0] Result_acc_170_nl;
  wire[19:0] nl_Result_acc_170_nl;
  wire[22:0] Result_acc_253_nl;
  wire[23:0] nl_Result_acc_253_nl;
  wire[17:0] MultLoop_acc_464_nl;
  wire[18:0] nl_MultLoop_acc_464_nl;
  wire[20:0] Result_acc_205_nl;
  wire[21:0] nl_Result_acc_205_nl;
  wire[17:0] Result_acc_204_nl;
  wire[18:0] nl_Result_acc_204_nl;
  wire[22:0] Result_acc_186_nl;
  wire[23:0] nl_Result_acc_186_nl;
  wire[19:0] Result_acc_185_nl;
  wire[20:0] nl_Result_acc_185_nl;
  wire[9:0] Result_acc_203_nl;
  wire[10:0] nl_Result_acc_203_nl;
  wire[16:0] MultLoop_acc_461_nl;
  wire[17:0] nl_MultLoop_acc_461_nl;
  wire[22:0] Result_acc_10_nl;
  wire[23:0] nl_Result_acc_10_nl;
  wire[14:0] Result_acc_206_nl;
  wire[15:0] nl_Result_acc_206_nl;
  wire[22:0] Result_acc_11_nl;
  wire[23:0] nl_Result_acc_11_nl;
  wire[21:0] Result_acc_174_nl;
  wire[23:0] nl_Result_acc_174_nl;
  wire[23:0] Result_acc_17_nl;
  wire[24:0] nl_Result_acc_17_nl;
  wire[22:0] Result_acc_179_nl;
  wire[24:0] nl_Result_acc_179_nl;
  wire[22:0] Result_acc_16_nl;
  wire[23:0] nl_Result_acc_16_nl;
  wire[20:0] Result_acc_176_nl;
  wire[21:0] nl_Result_acc_176_nl;
  wire[13:0] MultLoop_acc_458_nl;
  wire[14:0] nl_MultLoop_acc_458_nl;
  wire[22:0] Result_acc_8_nl;
  wire[23:0] nl_Result_acc_8_nl;
  wire[19:0] Result_acc_167_nl;
  wire[20:0] nl_Result_acc_167_nl;
  wire[13:0] Result_acc_208_nl;
  wire[14:0] nl_Result_acc_208_nl;
  wire[19:0] Result_acc_15_nl;
  wire[20:0] nl_Result_acc_15_nl;
  wire[17:0] Result_acc_168_nl;
  wire[18:0] nl_Result_acc_168_nl;
  wire[17:0] MultLoop_acc_1013_nl;
  wire[19:0] nl_MultLoop_acc_1013_nl;
  wire[17:0] MultLoop_acc_1011_nl;
  wire[18:0] nl_MultLoop_acc_1011_nl;
  wire[23:0] MultLoop_acc_311_nl;
  wire[24:0] nl_MultLoop_acc_311_nl;
  wire[22:0] MultLoop_acc_1005_nl;
  wire[23:0] nl_MultLoop_acc_1005_nl;
  wire[16:0] MultLoop_acc_1009_nl;
  wire[18:0] nl_MultLoop_acc_1009_nl;
  wire[21:0] MultLoop_acc_1394_nl;
  wire[22:0] nl_MultLoop_acc_1394_nl;
  wire[17:0] MultLoop_acc_75_nl;
  wire[18:0] nl_MultLoop_acc_75_nl;
  wire[13:0] MultLoop_acc_1006_nl;
  wire[14:0] nl_MultLoop_acc_1006_nl;
  wire[19:0] MultLoop_acc_1383_nl;
  wire[20:0] nl_MultLoop_acc_1383_nl;
  wire[23:0] MultLoop_acc_73_nl;
  wire[25:0] nl_MultLoop_acc_73_nl;
  wire[13:0] MultLoop_acc_1302_nl;
  wire[14:0] nl_MultLoop_acc_1302_nl;
  wire[17:0] MultLoop_acc_1305_nl;
  wire[18:0] nl_MultLoop_acc_1305_nl;
  wire[18:0] MultLoop_acc_1304_nl;
  wire[19:0] nl_MultLoop_acc_1304_nl;
  wire[17:0] MultLoop_acc_1012_nl;
  wire[18:0] nl_MultLoop_acc_1012_nl;
  wire[18:0] MultLoop_acc_1306_nl;
  wire[19:0] nl_MultLoop_acc_1306_nl;
  wire[24:0] MultLoop_acc_1001_nl;
  wire[25:0] nl_MultLoop_acc_1001_nl;
  wire[21:0] MultLoop_acc_1000_nl;
  wire[22:0] nl_MultLoop_acc_1000_nl;
  wire[19:0] MultLoop_acc_1308_nl;
  wire[20:0] nl_MultLoop_acc_1308_nl;
  wire[17:0] MultLoop_acc_1307_nl;
  wire[18:0] nl_MultLoop_acc_1307_nl;
  wire[17:0] MultLoop_acc_483_nl;
  wire[18:0] nl_MultLoop_acc_483_nl;
  wire[17:0] MultLoop_acc_481_nl;
  wire[18:0] nl_MultLoop_acc_481_nl;
  wire[17:0] MultLoop_acc_477_nl;
  wire[18:0] nl_MultLoop_acc_477_nl;
  wire[17:0] Result_acc_199_nl;
  wire[18:0] nl_Result_acc_199_nl;
  wire[18:0] Result_acc_250_nl;
  wire[19:0] nl_Result_acc_250_nl;
  wire[19:0] MultLoop_acc_1381_nl;
  wire[20:0] nl_MultLoop_acc_1381_nl;
  wire[18:0] MultLoop_acc_1298_nl;
  wire[19:0] nl_MultLoop_acc_1298_nl;
  wire[18:0] MultLoop_acc_1382_nl;
  wire[19:0] nl_MultLoop_acc_1382_nl;
  wire[17:0] MultLoop_acc_480_nl;
  wire[18:0] nl_MultLoop_acc_480_nl;
  wire[18:0] Result_acc_nl;
  wire[19:0] nl_Result_acc_nl;
  wire[23:0] Result_acc_194_nl;
  wire[24:0] nl_Result_acc_194_nl;
  wire[19:0] Result_acc_201_nl;
  wire[20:0] nl_Result_acc_201_nl;
  wire[17:0] Result_acc_200_nl;
  wire[18:0] nl_Result_acc_200_nl;
  wire[21:0] Result_acc_196_nl;
  wire[22:0] nl_Result_acc_196_nl;
  wire[17:0] MultLoop_acc_1301_nl;
  wire[18:0] nl_MultLoop_acc_1301_nl;
  wire[21:0] MultLoop_acc_470_nl;
  wire[22:0] nl_MultLoop_acc_470_nl;
  wire[17:0] MultLoop_acc_469_nl;
  wire[18:0] nl_MultLoop_acc_469_nl;
  wire[18:0] MultLoop_acc_1299_nl;
  wire[19:0] nl_MultLoop_acc_1299_nl;
  wire[21:0] MultLoop_acc_467_nl;
  wire[22:0] nl_MultLoop_acc_467_nl;
  wire[13:0] MultLoop_acc_278_nl;
  wire[14:0] nl_MultLoop_acc_278_nl;
  wire[25:0] MultLoop_acc_284_nl;
  wire[26:0] nl_MultLoop_acc_284_nl;
  wire[24:0] MultLoop_acc_472_nl;
  wire[26:0] nl_MultLoop_acc_472_nl;
  wire[22:0] Result_acc_2_nl;
  wire[23:0] nl_Result_acc_2_nl;
  wire[20:0] Result_acc_190_nl;
  wire[21:0] nl_Result_acc_190_nl;
  wire[17:0] Result_acc_189_nl;
  wire[18:0] nl_Result_acc_189_nl;
  wire[17:0] MultLoop_acc_989_nl;
  wire[18:0] nl_MultLoop_acc_989_nl;
  wire[17:0] MultLoop_acc_986_nl;
  wire[18:0] nl_MultLoop_acc_986_nl;
  wire[21:0] MultLoop_acc_1380_nl;
  wire[22:0] nl_MultLoop_acc_1380_nl;
  wire[15:0] MultLoop_acc_984_nl;
  wire[17:0] nl_MultLoop_acc_984_nl;
  wire[25:0] MultLoop_acc_82_nl;
  wire[26:0] nl_MultLoop_acc_82_nl;
  wire[21:0] MultLoop_acc_973_nl;
  wire[22:0] nl_MultLoop_acc_973_nl;
  wire[19:0] MultLoop_acc_972_nl;
  wire[20:0] nl_MultLoop_acc_972_nl;
  wire[23:0] MultLoop_acc_77_nl;
  wire[24:0] nl_MultLoop_acc_77_nl;
  wire[21:0] MultLoop_acc_966_nl;
  wire[22:0] nl_MultLoop_acc_966_nl;
  wire[21:0] MultLoop_acc_78_nl;
  wire[22:0] nl_MultLoop_acc_78_nl;
  wire[19:0] MultLoop_acc_964_nl;
  wire[20:0] nl_MultLoop_acc_964_nl;
  wire[14:0] MultLoop_acc_1297_nl;
  wire[15:0] nl_MultLoop_acc_1297_nl;
  wire[21:0] MultLoop_acc_86_nl;
  wire[22:0] nl_MultLoop_acc_86_nl;
  wire[18:0] MultLoop_acc_975_nl;
  wire[19:0] nl_MultLoop_acc_975_nl;
  wire[17:0] MultLoop_acc_1293_nl;
  wire[18:0] nl_MultLoop_acc_1293_nl;
  wire[21:0] MultLoop_acc_315_nl;
  wire[22:0] nl_MultLoop_acc_315_nl;
  wire[20:0] MultLoop_acc_970_nl;
  wire[21:0] nl_MultLoop_acc_970_nl;
  wire[17:0] MultLoop_acc_969_nl;
  wire[18:0] nl_MultLoop_acc_969_nl;
  wire[26:0] MultLoop_acc_83_nl;
  wire[27:0] nl_MultLoop_acc_83_nl;
  wire[21:0] MultLoop_acc_976_nl;
  wire[22:0] nl_MultLoop_acc_976_nl;
  wire[22:0] MultLoop_acc_79_nl;
  wire[24:0] nl_MultLoop_acc_79_nl;
  wire[14:0] MultLoop_acc_1295_nl;
  wire[15:0] nl_MultLoop_acc_1295_nl;
  wire[17:0] MultLoop_acc_510_nl;
  wire[19:0] nl_MultLoop_acc_510_nl;
  wire[18:0] MultLoop_acc_1287_nl;
  wire[19:0] nl_MultLoop_acc_1287_nl;
  wire[23:0] MultLoop_acc_496_nl;
  wire[25:0] nl_MultLoop_acc_496_nl;
  wire[16:0] MultLoop_242_MultLoop_acc_3_nl;
  wire[17:0] nl_MultLoop_242_MultLoop_acc_3_nl;
  wire[13:0] MultLoop_acc_501_nl;
  wire[14:0] nl_MultLoop_acc_501_nl;
  wire[20:0] MultLoop_acc_1290_nl;
  wire[21:0] nl_MultLoop_acc_1290_nl;
  wire[17:0] MultLoop_acc_1289_nl;
  wire[18:0] nl_MultLoop_acc_1289_nl;
  wire[21:0] MultLoop_acc_499_nl;
  wire[23:0] nl_MultLoop_acc_499_nl;
  wire[20:0] MultLoop_acc_270_nl;
  wire[21:0] nl_MultLoop_acc_270_nl;
  wire[16:0] MultLoop_acc_1291_nl;
  wire[17:0] nl_MultLoop_acc_1291_nl;
  wire[23:0] MultLoop_acc_1379_nl;
  wire[24:0] nl_MultLoop_acc_1379_nl;
  wire[17:0] MultLoop_acc_509_nl;
  wire[18:0] nl_MultLoop_acc_509_nl;
  wire[19:0] MultLoop_acc_269_nl;
  wire[20:0] nl_MultLoop_acc_269_nl;
  wire[18:0] MultLoop_acc_504_nl;
  wire[19:0] nl_MultLoop_acc_504_nl;
  wire[14:0] MultLoop_acc_1282_nl;
  wire[15:0] nl_MultLoop_acc_1282_nl;
  wire[16:0] MultLoop_acc_505_nl;
  wire[17:0] nl_MultLoop_acc_505_nl;
  wire[17:0] MultLoop_acc_1284_nl;
  wire[18:0] nl_MultLoop_acc_1284_nl;
  wire[18:0] MultLoop_acc_1393_nl;
  wire[19:0] nl_MultLoop_acc_1393_nl;
  wire[24:0] MultLoop_acc_271_nl;
  wire[25:0] nl_MultLoop_acc_271_nl;
  wire[21:0] MultLoop_acc_485_nl;
  wire[22:0] nl_MultLoop_acc_485_nl;
  wire[20:0] MultLoop_acc_365_nl;
  wire[21:0] nl_MultLoop_acc_365_nl;
  wire[18:0] MultLoop_acc_490_nl;
  wire[19:0] nl_MultLoop_acc_490_nl;
  wire[17:0] MultLoop_acc_1286_nl;
  wire[18:0] nl_MultLoop_acc_1286_nl;
  wire[19:0] MultLoop_acc_493_nl;
  wire[20:0] nl_MultLoop_acc_493_nl;
  wire[17:0] MultLoop_acc_492_nl;
  wire[18:0] nl_MultLoop_acc_492_nl;
  wire[17:0] MultLoop_acc_961_nl;
  wire[19:0] nl_MultLoop_acc_961_nl;
  wire[26:0] MultLoop_acc_95_nl;
  wire[27:0] nl_MultLoop_acc_95_nl;
  wire[10:0] MultLoop_acc_1278_nl;
  wire[11:0] nl_MultLoop_acc_1278_nl;
  wire[17:0] MultLoop_acc_1281_nl;
  wire[18:0] nl_MultLoop_acc_1281_nl;
  wire[18:0] MultLoop_acc_1280_nl;
  wire[19:0] nl_MultLoop_acc_1280_nl;
  wire[22:0] MultLoop_acc_947_nl;
  wire[24:0] nl_MultLoop_acc_947_nl;
  wire[9:0] MultLoop_acc_1279_nl;
  wire[10:0] nl_MultLoop_acc_1279_nl;
  wire[16:0] MultLoop_71_MultLoop_acc_3_nl;
  wire[17:0] nl_MultLoop_71_MultLoop_acc_3_nl;
  wire[17:0] MultLoop_acc_960_nl;
  wire[18:0] nl_MultLoop_acc_960_nl;
  wire[17:0] MultLoop_acc_956_nl;
  wire[18:0] nl_MultLoop_acc_956_nl;
  wire[18:0] MultLoop_acc_1377_nl;
  wire[19:0] nl_MultLoop_acc_1377_nl;
  wire[20:0] MultLoop_acc_317_nl;
  wire[21:0] nl_MultLoop_acc_317_nl;
  wire[23:0] MultLoop_acc_318_nl;
  wire[24:0] nl_MultLoop_acc_318_nl;
  wire[19:0] MultLoop_acc_951_nl;
  wire[20:0] nl_MultLoop_acc_951_nl;
  wire[17:0] MultLoop_acc_950_nl;
  wire[18:0] nl_MultLoop_acc_950_nl;
  wire[17:0] MultLoop_acc_959_nl;
  wire[18:0] nl_MultLoop_acc_959_nl;
  wire[17:0] MultLoop_acc_1274_nl;
  wire[18:0] nl_MultLoop_acc_1274_nl;
  wire[20:0] MultLoop_acc_954_nl;
  wire[22:0] nl_MultLoop_acc_954_nl;
  wire[16:0] MultLoop_acc_955_nl;
  wire[17:0] nl_MultLoop_acc_955_nl;
  wire[19:0] MultLoop_acc_93_nl;
  wire[20:0] nl_MultLoop_acc_93_nl;
  wire[18:0] MultLoop_acc_942_nl;
  wire[19:0] nl_MultLoop_acc_942_nl;
  wire[12:0] MultLoop_acc_1275_nl;
  wire[13:0] nl_MultLoop_acc_1275_nl;
  wire[17:0] MultLoop_acc_1277_nl;
  wire[18:0] nl_MultLoop_acc_1277_nl;
  wire[19:0] MultLoop_acc_1411_nl;
  wire[20:0] nl_MultLoop_acc_1411_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_13_nl;
  wire[19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_13_nl;
  wire[24:0] MultLoop_acc_260_nl;
  wire[25:0] nl_MultLoop_acc_260_nl;
  wire[23:0] MultLoop_acc_525_nl;
  wire[24:0] nl_MultLoop_acc_525_nl;
  wire[25:0] MultLoop_acc_263_nl;
  wire[26:0] nl_MultLoop_acc_263_nl;
  wire[23:0] MultLoop_acc_521_nl;
  wire[25:0] nl_MultLoop_acc_521_nl;
  wire[22:0] MultLoop_acc_1406_nl;
  wire[23:0] nl_MultLoop_acc_1406_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_12_nl;
  wire[18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_12_nl;
  wire[20:0] MultLoop_acc_1268_nl;
  wire[21:0] nl_MultLoop_acc_1268_nl;
  wire[17:0] MultLoop_acc_1267_nl;
  wire[18:0] nl_MultLoop_acc_1267_nl;
  wire[20:0] MultLoop_acc_526_nl;
  wire[21:0] nl_MultLoop_acc_526_nl;
  wire[16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_9_nl;
  wire[17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_9_nl;
  wire[15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_7_nl;
  wire[17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_7_nl;
  wire[21:0] MultLoop_acc_259_nl;
  wire[22:0] nl_MultLoop_acc_259_nl;
  wire[18:0] MultLoop_acc_513_nl;
  wire[19:0] nl_MultLoop_acc_513_nl;
  wire[12:0] MultLoop_acc_1269_nl;
  wire[13:0] nl_MultLoop_acc_1269_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_nor_nl;
  wire[23:0] MultLoop_acc_364_nl;
  wire[24:0] nl_MultLoop_acc_364_nl;
  wire[21:0] MultLoop_acc_515_nl;
  wire[22:0] nl_MultLoop_acc_515_nl;
  wire[17:0] MultLoop_acc_1271_nl;
  wire[18:0] nl_MultLoop_acc_1271_nl;
  wire[21:0] MultLoop_acc_519_nl;
  wire[22:0] nl_MultLoop_acc_519_nl;
  wire[12:0] MultLoop_acc_1270_nl;
  wire[13:0] nl_MultLoop_acc_1270_nl;
  wire[15:0] MultLoop_231_MultLoop_acc_3_nl;
  wire[16:0] nl_MultLoop_231_MultLoop_acc_3_nl;
  wire[20:0] MultLoop_acc_1376_nl;
  wire[21:0] nl_MultLoop_acc_1376_nl;
  wire[17:0] MultLoop_acc_935_nl;
  wire[19:0] nl_MultLoop_acc_935_nl;
  wire[25:0] MultLoop_acc_104_nl;
  wire[26:0] nl_MultLoop_acc_104_nl;
  wire[24:0] MultLoop_acc_925_nl;
  wire[26:0] nl_MultLoop_acc_925_nl;
  wire[14:0] MultLoop_acc_99_nl;
  wire[15:0] nl_MultLoop_acc_99_nl;
  wire[17:0] MultLoop_acc_1266_nl;
  wire[18:0] nl_MultLoop_acc_1266_nl;
  wire[18:0] MultLoop_acc_1392_nl;
  wire[19:0] nl_MultLoop_acc_1392_nl;
  wire[17:0] MultLoop_acc_934_nl;
  wire[18:0] nl_MultLoop_acc_934_nl;
  wire[25:0] MultLoop_acc_321_nl;
  wire[26:0] nl_MultLoop_acc_321_nl;
  wire[24:0] MultLoop_acc_928_nl;
  wire[25:0] nl_MultLoop_acc_928_nl;
  wire[21:0] MultLoop_acc_927_nl;
  wire[22:0] nl_MultLoop_acc_927_nl;
  wire[16:0] MultLoop_acc_931_nl;
  wire[17:0] nl_MultLoop_acc_931_nl;
  wire[22:0] MultLoop_acc_320_nl;
  wire[23:0] nl_MultLoop_acc_320_nl;
  wire[18:0] MultLoop_acc_918_nl;
  wire[19:0] nl_MultLoop_acc_918_nl;
  wire[24:0] MultLoop_acc_103_nl;
  wire[26:0] nl_MultLoop_acc_103_nl;
  wire[19:0] MultLoop_acc_919_nl;
  wire[20:0] nl_MultLoop_acc_919_nl;
  wire[18:0] MultLoop_acc_1264_nl;
  wire[19:0] nl_MultLoop_acc_1264_nl;
  wire[19:0] MultLoop_acc_922_nl;
  wire[20:0] nl_MultLoop_acc_922_nl;
  wire[24:0] MultLoop_acc_101_nl;
  wire[25:0] nl_MultLoop_acc_101_nl;
  wire[22:0] MultLoop_acc_921_nl;
  wire[23:0] nl_MultLoop_acc_921_nl;
  wire[19:0] MultLoop_acc_319_nl;
  wire[20:0] nl_MultLoop_acc_319_nl;
  wire[17:0] MultLoop_acc_914_nl;
  wire[18:0] nl_MultLoop_acc_914_nl;
  wire[17:0] MultLoop_acc_553_nl;
  wire[18:0] nl_MultLoop_acc_553_nl;
  wire[17:0] MultLoop_acc_551_nl;
  wire[18:0] nl_MultLoop_acc_551_nl;
  wire[20:0] MultLoop_acc_360_nl;
  wire[21:0] nl_MultLoop_acc_360_nl;
  wire[17:0] MultLoop_acc_542_nl;
  wire[18:0] nl_MultLoop_acc_542_nl;
  wire[18:0] MultLoop_acc_1256_nl;
  wire[19:0] nl_MultLoop_acc_1256_nl;
  wire[21:0] MultLoop_acc_544_nl;
  wire[22:0] nl_MultLoop_acc_544_nl;
  wire[17:0] MultLoop_acc_550_nl;
  wire[19:0] nl_MultLoop_acc_550_nl;
  wire[22:0] MultLoop_acc_254_nl;
  wire[23:0] nl_MultLoop_acc_254_nl;
  wire[21:0] MultLoop_acc_529_nl;
  wire[22:0] nl_MultLoop_acc_529_nl;
  wire[17:0] MultLoop_acc_1258_nl;
  wire[18:0] nl_MultLoop_acc_1258_nl;
  wire[22:0] MultLoop_acc_532_nl;
  wire[23:0] nl_MultLoop_acc_532_nl;
  wire[19:0] MultLoop_acc_531_nl;
  wire[20:0] nl_MultLoop_acc_531_nl;
  wire[18:0] MultLoop_acc_362_nl;
  wire[19:0] nl_MultLoop_acc_362_nl;
  wire[12:0] MultLoop_acc_545_nl;
  wire[13:0] nl_MultLoop_acc_545_nl;
  wire[21:0] MultLoop_acc_253_nl;
  wire[22:0] nl_MultLoop_acc_253_nl;
  wire[15:0] MultLoop_acc_1259_nl;
  wire[16:0] nl_MultLoop_acc_1259_nl;
  wire[21:0] MultLoop_acc_363_nl;
  wire[22:0] nl_MultLoop_acc_363_nl;
  wire[20:0] MultLoop_acc_534_nl;
  wire[21:0] nl_MultLoop_acc_534_nl;
  wire[17:0] MultLoop_acc_533_nl;
  wire[18:0] nl_MultLoop_acc_533_nl;
  wire[17:0] MultLoop_acc_1262_nl;
  wire[18:0] nl_MultLoop_acc_1262_nl;
  wire[18:0] MultLoop_acc_1261_nl;
  wire[19:0] nl_MultLoop_acc_1261_nl;
  wire[18:0] MultLoop_acc_1410_nl;
  wire[19:0] nl_MultLoop_acc_1410_nl;
  wire[19:0] MultLoop_acc_1263_nl;
  wire[20:0] nl_MultLoop_acc_1263_nl;
  wire[20:0] MultLoop_acc_1375_nl;
  wire[21:0] nl_MultLoop_acc_1375_nl;
  wire[22:0] MultLoop_acc_255_nl;
  wire[23:0] nl_MultLoop_acc_255_nl;
  wire[17:0] MultLoop_acc_913_nl;
  wire[18:0] nl_MultLoop_acc_913_nl;
  wire[17:0] MultLoop_acc_911_nl;
  wire[18:0] nl_MultLoop_acc_911_nl;
  wire[16:0] MultLoop_acc_1248_nl;
  wire[17:0] nl_MultLoop_acc_1248_nl;
  wire[20:0] MultLoop_acc_1251_nl;
  wire[21:0] nl_MultLoop_acc_1251_nl;
  wire[17:0] MultLoop_acc_1250_nl;
  wire[18:0] nl_MultLoop_acc_1250_nl;
  wire[20:0] MultLoop_acc_903_nl;
  wire[21:0] nl_MultLoop_acc_903_nl;
  wire[17:0] MultLoop_acc_910_nl;
  wire[18:0] nl_MultLoop_acc_910_nl;
  wire[15:0] MultLoop_acc_907_nl;
  wire[16:0] nl_MultLoop_acc_907_nl;
  wire[14:0] MultLoop_acc_905_nl;
  wire[15:0] nl_MultLoop_acc_905_nl;
  wire[17:0] MultLoop_acc_111_nl;
  wire[18:0] nl_MultLoop_acc_111_nl;
  wire[19:0] MultLoop_acc_1253_nl;
  wire[20:0] nl_MultLoop_acc_1253_nl;
  wire[17:0] MultLoop_acc_1252_nl;
  wire[18:0] nl_MultLoop_acc_1252_nl;
  wire[17:0] MultLoop_acc_912_nl;
  wire[19:0] nl_MultLoop_acc_912_nl;
  wire[16:0] MultLoop_acc_908_nl;
  wire[17:0] nl_MultLoop_acc_908_nl;
  wire[15:0] MultLoop_acc_906_nl;
  wire[16:0] nl_MultLoop_acc_906_nl;
  wire[21:0] MultLoop_acc_117_nl;
  wire[22:0] nl_MultLoop_acc_117_nl;
  wire[22:0] MultLoop_acc_110_nl;
  wire[23:0] nl_MultLoop_acc_110_nl;
  wire[18:0] MultLoop_acc_891_nl;
  wire[19:0] nl_MultLoop_acc_891_nl;
  wire[24:0] MultLoop_acc_324_nl;
  wire[25:0] nl_MultLoop_acc_324_nl;
  wire[22:0] MultLoop_acc_897_nl;
  wire[23:0] nl_MultLoop_acc_897_nl;
  wire[20:0] MultLoop_acc_896_nl;
  wire[21:0] nl_MultLoop_acc_896_nl;
  wire[17:0] MultLoop_acc_577_nl;
  wire[18:0] nl_MultLoop_acc_577_nl;
  wire[17:0] MultLoop_acc_575_nl;
  wire[18:0] nl_MultLoop_acc_575_nl;
  wire[20:0] MultLoop_acc_1391_nl;
  wire[21:0] nl_MultLoop_acc_1391_nl;
  wire[22:0] MultLoop_acc_359_nl;
  wire[23:0] nl_MultLoop_acc_359_nl;
  wire[20:0] MultLoop_acc_568_nl;
  wire[21:0] nl_MultLoop_acc_568_nl;
  wire[17:0] MultLoop_acc_567_nl;
  wire[18:0] nl_MultLoop_acc_567_nl;
  wire[17:0] MultLoop_acc_574_nl;
  wire[20:0] nl_MultLoop_acc_574_nl;
  wire[18:0] MultLoop_acc_1371_nl;
  wire[19:0] nl_MultLoop_acc_1371_nl;
  wire[19:0] MultLoop_acc_1372_nl;
  wire[20:0] nl_MultLoop_acc_1372_nl;
  wire[22:0] MultLoop_acc_356_nl;
  wire[23:0] nl_MultLoop_acc_356_nl;
  wire[14:0] MultLoop_acc_569_nl;
  wire[15:0] nl_MultLoop_acc_569_nl;
  wire[19:0] MultLoop_acc_1370_nl;
  wire[20:0] nl_MultLoop_acc_1370_nl;
  wire[27:0] MultLoop_acc_240_nl;
  wire[29:0] nl_MultLoop_acc_240_nl;
  wire[23:0] MultLoop_acc_358_nl;
  wire[24:0] nl_MultLoop_acc_358_nl;
  wire[21:0] MultLoop_acc_559_nl;
  wire[22:0] nl_MultLoop_acc_559_nl;
  wire[17:0] MultLoop_acc_558_nl;
  wire[18:0] nl_MultLoop_acc_558_nl;
  wire[18:0] MultLoop_acc_1245_nl;
  wire[19:0] nl_MultLoop_acc_1245_nl;
  wire[20:0] MultLoop_acc_1373_nl;
  wire[21:0] nl_MultLoop_acc_1373_nl;
  wire[17:0] MultLoop_acc_889_nl;
  wire[18:0] nl_MultLoop_acc_889_nl;
  wire[17:0] MultLoop_acc_887_nl;
  wire[18:0] nl_MultLoop_acc_887_nl;
  wire[18:0] MultLoop_acc_1237_nl;
  wire[19:0] nl_MultLoop_acc_1237_nl;
  wire[20:0] MultLoop_acc_1368_nl;
  wire[21:0] nl_MultLoop_acc_1368_nl;
  wire[23:0] MultLoop_acc_127_nl;
  wire[24:0] nl_MultLoop_acc_127_nl;
  wire[19:0] MultLoop_acc_880_nl;
  wire[20:0] nl_MultLoop_acc_880_nl;
  wire[17:0] MultLoop_acc_886_nl;
  wire[18:0] nl_MultLoop_acc_886_nl;
  wire[18:0] MultLoop_acc_1238_nl;
  wire[19:0] nl_MultLoop_acc_1238_nl;
  wire[21:0] MultLoop_acc_881_nl;
  wire[22:0] nl_MultLoop_acc_881_nl;
  wire[16:0] MultLoop_acc_884_nl;
  wire[18:0] nl_MultLoop_acc_884_nl;
  wire[14:0] MultLoop_101_MultLoop_acc_3_nl;
  wire[15:0] nl_MultLoop_101_MultLoop_acc_3_nl;
  wire[20:0] MultLoop_acc_120_nl;
  wire[21:0] nl_MultLoop_acc_120_nl;
  wire[18:0] MultLoop_acc_867_nl;
  wire[19:0] nl_MultLoop_acc_867_nl;
  wire[17:0] MultLoop_acc_124_nl;
  wire[18:0] nl_MultLoop_acc_124_nl;
  wire[17:0] MultLoop_acc_888_nl;
  wire[18:0] nl_MultLoop_acc_888_nl;
  wire[17:0] MultLoop_acc_885_nl;
  wire[18:0] nl_MultLoop_acc_885_nl;
  wire[17:0] MultLoop_acc_1241_nl;
  wire[18:0] nl_MultLoop_acc_1241_nl;
  wire[23:0] MultLoop_acc_871_nl;
  wire[24:0] nl_MultLoop_acc_871_nl;
  wire[21:0] MultLoop_acc_870_nl;
  wire[22:0] nl_MultLoop_acc_870_nl;
  wire[19:0] MultLoop_acc_869_nl;
  wire[20:0] nl_MultLoop_acc_869_nl;
  wire[9:0] MultLoop_acc_1240_nl;
  wire[10:0] nl_MultLoop_acc_1240_nl;
  wire[17:0] MultLoop_acc_1243_nl;
  wire[18:0] nl_MultLoop_acc_1243_nl;
  wire[23:0] MultLoop_acc_874_nl;
  wire[25:0] nl_MultLoop_acc_874_nl;
  wire[18:0] MultLoop_acc_1244_nl;
  wire[19:0] nl_MultLoop_acc_1244_nl;
  wire[18:0] MultLoop_acc_1369_nl;
  wire[19:0] nl_MultLoop_acc_1369_nl;
  wire[17:0] MultLoop_acc_603_nl;
  wire[19:0] nl_MultLoop_acc_603_nl;
  wire[17:0] MultLoop_acc_1233_nl;
  wire[18:0] nl_MultLoop_acc_1233_nl;
  wire[24:0] MultLoop_acc_587_nl;
  wire[26:0] nl_MultLoop_acc_587_nl;
  wire[17:0] MultLoop_acc_1235_nl;
  wire[18:0] nl_MultLoop_acc_1235_nl;
  wire[24:0] MultLoop_acc_591_nl;
  wire[26:0] nl_MultLoop_acc_591_nl;
  wire[16:0] MultLoop_202_MultLoop_acc_3_nl;
  wire[17:0] nl_MultLoop_202_MultLoop_acc_3_nl;
  wire[15:0] MultLoop_acc_595_nl;
  wire[16:0] nl_MultLoop_acc_595_nl;
  wire[23:0] MultLoop_acc_229_nl;
  wire[25:0] nl_MultLoop_acc_229_nl;
  wire[13:0] MultLoop_acc_1236_nl;
  wire[14:0] nl_MultLoop_acc_1236_nl;
  wire[18:0] MultLoop_acc_1407_nl;
  wire[19:0] nl_MultLoop_acc_1407_nl;
  wire[17:0] MultLoop_acc_602_nl;
  wire[18:0] nl_MultLoop_acc_602_nl;
  wire[18:0] MultLoop_acc_1231_nl;
  wire[19:0] nl_MultLoop_acc_1231_nl;
  wire[18:0] MultLoop_acc_1367_nl;
  wire[19:0] nl_MultLoop_acc_1367_nl;
  wire[16:0] MultLoop_acc_598_nl;
  wire[17:0] nl_MultLoop_acc_598_nl;
  wire[25:0] MultLoop_acc_232_nl;
  wire[26:0] nl_MultLoop_acc_232_nl;
  wire[23:0] MultLoop_acc_579_nl;
  wire[24:0] nl_MultLoop_acc_579_nl;
  wire[18:0] MultLoop_acc_1409_nl;
  wire[19:0] nl_MultLoop_acc_1409_nl;
  wire[20:0] MultLoop_acc_1389_nl;
  wire[21:0] nl_MultLoop_acc_1389_nl;
  wire[17:0] MultLoop_acc_864_nl;
  wire[18:0] nl_MultLoop_acc_864_nl;
  wire[17:0] MultLoop_acc_862_nl;
  wire[18:0] nl_MultLoop_acc_862_nl;
  wire[17:0] MultLoop_acc_858_nl;
  wire[18:0] nl_MultLoop_acc_858_nl;
  wire[22:0] MultLoop_acc_327_nl;
  wire[23:0] nl_MultLoop_acc_327_nl;
  wire[19:0] MultLoop_acc_836_nl;
  wire[21:0] nl_MultLoop_acc_836_nl;
  wire[12:0] MultLoop_acc_1222_nl;
  wire[13:0] nl_MultLoop_acc_1222_nl;
  wire[22:0] MultLoop_acc_328_nl;
  wire[23:0] nl_MultLoop_acc_328_nl;
  wire[19:0] MultLoop_acc_838_nl;
  wire[20:0] nl_MultLoop_acc_838_nl;
  wire[17:0] MultLoop_acc_837_nl;
  wire[18:0] nl_MultLoop_acc_837_nl;
  wire[19:0] MultLoop_acc_1223_nl;
  wire[20:0] nl_MultLoop_acc_1223_nl;
  wire[23:0] MultLoop_acc_1366_nl;
  wire[24:0] nl_MultLoop_acc_1366_nl;
  wire[17:0] MultLoop_acc_861_nl;
  wire[18:0] nl_MultLoop_acc_861_nl;
  wire[22:0] MultLoop_acc_133_nl;
  wire[23:0] nl_MultLoop_acc_133_nl;
  wire[20:0] MultLoop_acc_843_nl;
  wire[21:0] nl_MultLoop_acc_843_nl;
  wire[26:0] MultLoop_acc_134_nl;
  wire[27:0] nl_MultLoop_acc_134_nl;
  wire[21:0] MultLoop_acc_846_nl;
  wire[22:0] nl_MultLoop_acc_846_nl;
  wire[19:0] MultLoop_acc_845_nl;
  wire[20:0] nl_MultLoop_acc_845_nl;
  wire[17:0] MultLoop_acc_863_nl;
  wire[18:0] nl_MultLoop_acc_863_nl;
  wire[17:0] MultLoop_acc_860_nl;
  wire[18:0] nl_MultLoop_acc_860_nl;
  wire[24:0] MultLoop_acc_329_nl;
  wire[25:0] nl_MultLoop_acc_329_nl;
  wire[21:0] MultLoop_acc_849_nl;
  wire[23:0] nl_MultLoop_acc_849_nl;
  wire[19:0] MultLoop_acc_1227_nl;
  wire[20:0] nl_MultLoop_acc_1227_nl;
  wire[26:0] MultLoop_acc_853_nl;
  wire[28:0] nl_MultLoop_acc_853_nl;
  wire[17:0] MultLoop_acc_859_nl;
  wire[19:0] nl_MultLoop_acc_859_nl;
  wire[24:0] MultLoop_acc_140_nl;
  wire[25:0] nl_MultLoop_acc_140_nl;
  wire[21:0] MultLoop_acc_855_nl;
  wire[22:0] nl_MultLoop_acc_855_nl;
  wire[11:0] MultLoop_acc_1228_nl;
  wire[12:0] nl_MultLoop_acc_1228_nl;
  wire[22:0] MultLoop_acc_330_nl;
  wire[23:0] nl_MultLoop_acc_330_nl;
  wire[21:0] MultLoop_acc_833_nl;
  wire[22:0] nl_MultLoop_acc_833_nl;
  wire[17:0] MultLoop_acc_832_nl;
  wire[18:0] nl_MultLoop_acc_832_nl;
  wire[9:0] MultLoop_acc_1230_nl;
  wire[10:0] nl_MultLoop_acc_1230_nl;
  wire[17:0] MultLoop_acc_631_nl;
  wire[18:0] nl_MultLoop_acc_631_nl;
  wire[17:0] MultLoop_acc_629_nl;
  wire[18:0] nl_MultLoop_acc_629_nl;
  wire[18:0] MultLoop_acc_1363_nl;
  wire[19:0] nl_MultLoop_acc_1363_nl;
  wire[24:0] MultLoop_acc_352_nl;
  wire[25:0] nl_MultLoop_acc_352_nl;
  wire[21:0] MultLoop_acc_622_nl;
  wire[22:0] nl_MultLoop_acc_622_nl;
  wire[17:0] MultLoop_acc_628_nl;
  wire[18:0] nl_MultLoop_acc_628_nl;
  wire[18:0] MultLoop_acc_1364_nl;
  wire[19:0] nl_MultLoop_acc_1364_nl;
  wire[16:0] MultLoop_acc_625_nl;
  wire[17:0] nl_MultLoop_acc_625_nl;
  wire[25:0] MultLoop_acc_220_nl;
  wire[26:0] nl_MultLoop_acc_220_nl;
  wire[22:0] MultLoop_acc_619_nl;
  wire[23:0] nl_MultLoop_acc_619_nl;
  wire[19:0] MultLoop_acc_618_nl;
  wire[20:0] nl_MultLoop_acc_618_nl;
  wire[25:0] MultLoop_acc_221_nl;
  wire[26:0] nl_MultLoop_acc_221_nl;
  wire[24:0] MultLoop_acc_605_nl;
  wire[25:0] nl_MultLoop_acc_605_nl;
  wire[24:0] MultLoop_acc_225_nl;
  wire[26:0] nl_MultLoop_acc_225_nl;
  wire[15:0] MultLoop_191_MultLoop_acc_3_nl;
  wire[16:0] nl_MultLoop_191_MultLoop_acc_3_nl;
  wire[18:0] MultLoop_acc_1365_nl;
  wire[19:0] nl_MultLoop_acc_1365_nl;
  wire[19:0] MultLoop_acc_1218_nl;
  wire[20:0] nl_MultLoop_acc_1218_nl;
  wire[17:0] MultLoop_acc_1217_nl;
  wire[18:0] nl_MultLoop_acc_1217_nl;
  wire[21:0] MultLoop_acc_608_nl;
  wire[23:0] nl_MultLoop_acc_608_nl;
  wire[17:0] MultLoop_acc_1221_nl;
  wire[18:0] nl_MultLoop_acc_1221_nl;
  wire[21:0] MultLoop_acc_613_nl;
  wire[22:0] nl_MultLoop_acc_613_nl;
  wire[12:0] MultLoop_acc_1220_nl;
  wire[13:0] nl_MultLoop_acc_1220_nl;
  wire[24:0] MultLoop_acc_350_nl;
  wire[25:0] nl_MultLoop_acc_350_nl;
  wire[22:0] MultLoop_acc_616_nl;
  wire[23:0] nl_MultLoop_acc_616_nl;
  wire[20:0] MultLoop_acc_615_nl;
  wire[21:0] nl_MultLoop_acc_615_nl;
  wire[17:0] MultLoop_acc_614_nl;
  wire[18:0] nl_MultLoop_acc_614_nl;
  wire[17:0] MultLoop_acc_830_nl;
  wire[20:0] nl_MultLoop_acc_830_nl;
  wire[19:0] MultLoop_acc_1362_nl;
  wire[20:0] nl_MultLoop_acc_1362_nl;
  wire[21:0] MultLoop_acc_331_nl;
  wire[22:0] nl_MultLoop_acc_331_nl;
  wire[19:0] MultLoop_acc_813_nl;
  wire[20:0] nl_MultLoop_acc_813_nl;
  wire[13:0] MultLoop_acc_822_nl;
  wire[14:0] nl_MultLoop_acc_822_nl;
  wire[21:0] MultLoop_acc_332_nl;
  wire[22:0] nl_MultLoop_acc_332_nl;
  wire[17:0] MultLoop_acc_804_nl;
  wire[18:0] nl_MultLoop_acc_804_nl;
  wire[13:0] MultLoop_acc_1212_nl;
  wire[14:0] nl_MultLoop_acc_1212_nl;
  wire[22:0] MultLoop_acc_334_nl;
  wire[23:0] nl_MultLoop_acc_334_nl;
  wire[17:0] MultLoop_acc_807_nl;
  wire[18:0] nl_MultLoop_acc_807_nl;
  wire[11:0] MultLoop_acc_1210_nl;
  wire[12:0] nl_MultLoop_acc_1210_nl;
  wire[18:0] MultLoop_acc_1360_nl;
  wire[19:0] nl_MultLoop_acc_1360_nl;
  wire[21:0] MultLoop_acc_1361_nl;
  wire[22:0] nl_MultLoop_acc_1361_nl;
  wire[19:0] MultLoop_acc_143_nl;
  wire[20:0] nl_MultLoop_acc_143_nl;
  wire[18:0] MultLoop_acc_811_nl;
  wire[19:0] nl_MultLoop_acc_811_nl;
  wire[17:0] MultLoop_acc_829_nl;
  wire[18:0] nl_MultLoop_acc_829_nl;
  wire[17:0] MultLoop_acc_1214_nl;
  wire[18:0] nl_MultLoop_acc_1214_nl;
  wire[23:0] MultLoop_acc_818_nl;
  wire[25:0] nl_MultLoop_acc_818_nl;
  wire[17:0] MultLoop_acc_816_nl;
  wire[18:0] nl_MultLoop_acc_816_nl;
  wire[17:0] MultLoop_acc_1215_nl;
  wire[18:0] nl_MultLoop_acc_1215_nl;
  wire[18:0] MultLoop_acc_1408_nl;
  wire[19:0] nl_MultLoop_acc_1408_nl;
  wire[17:0] MultLoop_acc_659_nl;
  wire[19:0] nl_MultLoop_acc_659_nl;
  wire[17:0] MultLoop_acc_657_nl;
  wire[18:0] nl_MultLoop_acc_657_nl;
  wire[22:0] MultLoop_acc_208_nl;
  wire[23:0] nl_MultLoop_acc_208_nl;
  wire[19:0] MultLoop_acc_643_nl;
  wire[20:0] nl_MultLoop_acc_643_nl;
  wire[27:0] MultLoop_acc_209_nl;
  wire[29:0] nl_MultLoop_acc_209_nl;
  wire[17:0] MultLoop_acc_1206_nl;
  wire[18:0] nl_MultLoop_acc_1206_nl;
  wire[23:0] MultLoop_acc_649_nl;
  wire[24:0] nl_MultLoop_acc_649_nl;
  wire[19:0] MultLoop_acc_648_nl;
  wire[20:0] nl_MultLoop_acc_648_nl;
  wire[17:0] MultLoop_acc_647_nl;
  wire[18:0] nl_MultLoop_acc_647_nl;
  wire[9:0] MultLoop_acc_1205_nl;
  wire[10:0] nl_MultLoop_acc_1205_nl;
  wire[23:0] MultLoop_acc_349_nl;
  wire[24:0] nl_MultLoop_acc_349_nl;
  wire[20:0] MultLoop_acc_651_nl;
  wire[21:0] nl_MultLoop_acc_651_nl;
  wire[17:0] MultLoop_acc_658_nl;
  wire[20:0] nl_MultLoop_acc_658_nl;
  wire[25:0] MultLoop_acc_211_nl;
  wire[26:0] nl_MultLoop_acc_211_nl;
  wire[22:0] MultLoop_acc_640_nl;
  wire[23:0] nl_MultLoop_acc_640_nl;
  wire[20:0] MultLoop_acc_639_nl;
  wire[21:0] nl_MultLoop_acc_639_nl;
  wire[15:0] MultLoop_acc_205_nl;
  wire[16:0] nl_MultLoop_acc_205_nl;
  wire[21:0] MultLoop_acc_215_nl;
  wire[22:0] nl_MultLoop_acc_215_nl;
  wire[19:0] MultLoop_acc_635_nl;
  wire[20:0] nl_MultLoop_acc_635_nl;
  wire[22:0] MultLoop_acc_207_nl;
  wire[23:0] nl_MultLoop_acc_207_nl;
  wire[18:0] MultLoop_acc_637_nl;
  wire[19:0] nl_MultLoop_acc_637_nl;
  wire[11:0] MultLoop_acc_1207_nl;
  wire[12:0] nl_MultLoop_acc_1207_nl;
  wire[24:0] MultLoop_acc_214_nl;
  wire[25:0] nl_MultLoop_acc_214_nl;
  wire[20:0] MultLoop_acc_632_nl;
  wire[21:0] nl_MultLoop_acc_632_nl;
  wire[17:0] MultLoop_acc_801_nl;
  wire[18:0] nl_MultLoop_acc_801_nl;
  wire[16:0] MultLoop_acc_1199_nl;
  wire[17:0] nl_MultLoop_acc_1199_nl;
  wire[16:0] MultLoop_acc_798_nl;
  wire[18:0] nl_MultLoop_acc_798_nl;
  wire[19:0] MultLoop_acc_1202_nl;
  wire[20:0] nl_MultLoop_acc_1202_nl;
  wire[17:0] MultLoop_acc_1201_nl;
  wire[18:0] nl_MultLoop_acc_1201_nl;
  wire[22:0] MultLoop_acc_158_nl;
  wire[24:0] nl_MultLoop_acc_158_nl;
  wire[14:0] MultLoop_acc_1200_nl;
  wire[15:0] nl_MultLoop_acc_1200_nl;
  wire[17:0] MultLoop_acc_1192_nl;
  wire[18:0] nl_MultLoop_acc_1192_nl;
  wire[18:0] MultLoop_acc_1387_nl;
  wire[19:0] nl_MultLoop_acc_1387_nl;
  wire[25:0] MultLoop_acc_155_nl;
  wire[27:0] nl_MultLoop_acc_155_nl;
  wire[18:0] MultLoop_acc_1194_nl;
  wire[19:0] nl_MultLoop_acc_1194_nl;
  wire[18:0] MultLoop_acc_1358_nl;
  wire[19:0] nl_MultLoop_acc_1358_nl;
  wire[17:0] MultLoop_acc_1196_nl;
  wire[18:0] nl_MultLoop_acc_1196_nl;
  wire[24:0] MultLoop_acc_791_nl;
  wire[25:0] nl_MultLoop_acc_791_nl;
  wire[21:0] MultLoop_acc_790_nl;
  wire[22:0] nl_MultLoop_acc_790_nl;
  wire[15:0] MultLoop_131_MultLoop_acc_3_nl;
  wire[16:0] nl_MultLoop_131_MultLoop_acc_3_nl;
  wire[19:0] MultLoop_acc_152_nl;
  wire[20:0] nl_MultLoop_acc_152_nl;
  wire[19:0] MultLoop_acc_335_nl;
  wire[20:0] nl_MultLoop_acc_335_nl;
  wire[17:0] MultLoop_acc_785_nl;
  wire[18:0] nl_MultLoop_acc_785_nl;
  wire[17:0] MultLoop_acc_687_nl;
  wire[19:0] nl_MultLoop_acc_687_nl;
  wire[18:0] MultLoop_acc_1181_nl;
  wire[19:0] nl_MultLoop_acc_1181_nl;
  wire[21:0] MultLoop_acc_669_nl;
  wire[22:0] nl_MultLoop_acc_669_nl;
  wire[17:0] MultLoop_acc_1183_nl;
  wire[18:0] nl_MultLoop_acc_1183_nl;
  wire[24:0] MultLoop_acc_674_nl;
  wire[25:0] nl_MultLoop_acc_674_nl;
  wire[21:0] MultLoop_acc_673_nl;
  wire[23:0] nl_MultLoop_acc_673_nl;
  wire[17:0] MultLoop_acc_671_nl;
  wire[18:0] nl_MultLoop_acc_671_nl;
  wire[8:0] MultLoop_acc_1182_nl;
  wire[9:0] nl_MultLoop_acc_1182_nl;
  wire[19:0] MultLoop_acc_1184_nl;
  wire[20:0] nl_MultLoop_acc_1184_nl;
  wire[26:0] MultLoop_acc_677_nl;
  wire[28:0] nl_MultLoop_acc_677_nl;
  wire[18:0] MultLoop_acc_1185_nl;
  wire[19:0] nl_MultLoop_acc_1185_nl;
  wire[18:0] MultLoop_acc_1356_nl;
  wire[19:0] nl_MultLoop_acc_1356_nl;
  wire[17:0] MultLoop_acc_686_nl;
  wire[18:0] nl_MultLoop_acc_686_nl;
  wire[17:0] MultLoop_acc_683_nl;
  wire[19:0] nl_MultLoop_acc_683_nl;
  wire[16:0] MultLoop_acc_682_nl;
  wire[17:0] nl_MultLoop_acc_682_nl;
  wire[17:0] MultLoop_acc_1187_nl;
  wire[18:0] nl_MultLoop_acc_1187_nl;
  wire[24:0] MultLoop_acc_664_nl;
  wire[25:0] nl_MultLoop_acc_664_nl;
  wire[21:0] MultLoop_acc_663_nl;
  wire[22:0] nl_MultLoop_acc_663_nl;
  wire[15:0] MultLoop_acc_680_nl;
  wire[16:0] nl_MultLoop_acc_680_nl;
  wire[14:0] MultLoop_171_MultLoop_acc_3_nl;
  wire[15:0] nl_MultLoop_171_MultLoop_acc_3_nl;
  wire[17:0] MultLoop_acc_194_nl;
  wire[18:0] nl_MultLoop_acc_194_nl;
  wire[21:0] MultLoop_acc_1357_nl;
  wire[22:0] nl_MultLoop_acc_1357_nl;
  wire[20:0] MultLoop_acc_346_nl;
  wire[21:0] nl_MultLoop_acc_346_nl;
  wire[17:0] MultLoop_acc_661_nl;
  wire[18:0] nl_MultLoop_acc_661_nl;
  wire[20:0] MultLoop_acc_1190_nl;
  wire[21:0] nl_MultLoop_acc_1190_nl;
  wire[17:0] MultLoop_acc_1189_nl;
  wire[18:0] nl_MultLoop_acc_1189_nl;
  wire[22:0] MultLoop_acc_667_nl;
  wire[24:0] nl_MultLoop_acc_667_nl;
  wire[17:0] MultLoop_acc_774_nl;
  wire[18:0] nl_MultLoop_acc_774_nl;
  wire[17:0] MultLoop_acc_772_nl;
  wire[18:0] nl_MultLoop_acc_772_nl;
  wire[19:0] MultLoop_acc_1173_nl;
  wire[20:0] nl_MultLoop_acc_1173_nl;
  wire[20:0] MultLoop_acc_1352_nl;
  wire[21:0] nl_MultLoop_acc_1352_nl;
  wire[17:0] MultLoop_acc_1172_nl;
  wire[18:0] nl_MultLoop_acc_1172_nl;
  wire[17:0] MultLoop_acc_1175_nl;
  wire[18:0] nl_MultLoop_acc_1175_nl;
  wire[24:0] MultLoop_acc_765_nl;
  wire[25:0] nl_MultLoop_acc_765_nl;
  wire[21:0] MultLoop_acc_764_nl;
  wire[22:0] nl_MultLoop_acc_764_nl;
  wire[17:0] MultLoop_acc_771_nl;
  wire[18:0] nl_MultLoop_acc_771_nl;
  wire[24:0] MultLoop_acc_339_nl;
  wire[25:0] nl_MultLoop_acc_339_nl;
  wire[22:0] MultLoop_acc_750_nl;
  wire[23:0] nl_MultLoop_acc_750_nl;
  wire[19:0] MultLoop_acc_749_nl;
  wire[21:0] nl_MultLoop_acc_749_nl;
  wire[18:0] MultLoop_acc_1353_nl;
  wire[19:0] nl_MultLoop_acc_1353_nl;
  wire[24:0] MultLoop_acc_337_nl;
  wire[25:0] nl_MultLoop_acc_337_nl;
  wire[21:0] MultLoop_acc_754_nl;
  wire[22:0] nl_MultLoop_acc_754_nl;
  wire[21:0] MultLoop_acc_165_nl;
  wire[22:0] nl_MultLoop_acc_165_nl;
  wire[19:0] MultLoop_acc_757_nl;
  wire[20:0] nl_MultLoop_acc_757_nl;
  wire[17:0] MultLoop_acc_756_nl;
  wire[18:0] nl_MultLoop_acc_756_nl;
  wire[19:0] MultLoop_acc_336_nl;
  wire[20:0] nl_MultLoop_acc_336_nl;
  wire[17:0] MultLoop_acc_758_nl;
  wire[18:0] nl_MultLoop_acc_758_nl;
  wire[15:0] MultLoop_acc_768_nl;
  wire[16:0] nl_MultLoop_acc_768_nl;
  wire[18:0] MultLoop_acc_1179_nl;
  wire[19:0] nl_MultLoop_acc_1179_nl;
  wire[13:0] MultLoop_acc_767_nl;
  wire[14:0] nl_MultLoop_acc_767_nl;
  wire[20:0] MultLoop_acc_1355_nl;
  wire[21:0] nl_MultLoop_acc_1355_nl;
  wire[8:0] MultLoop_acc_1180_nl;
  wire[9:0] nl_MultLoop_acc_1180_nl;
  wire[17:0] MultLoop_acc_712_nl;
  wire[19:0] nl_MultLoop_acc_712_nl;
  wire[18:0] MultLoop_acc_1165_nl;
  wire[19:0] nl_MultLoop_acc_1165_nl;
  wire[24:0] MultLoop_acc_696_nl;
  wire[26:0] nl_MultLoop_acc_696_nl;
  wire[18:0] MultLoop_acc_1166_nl;
  wire[19:0] nl_MultLoop_acc_1166_nl;
  wire[21:0] MultLoop_acc_698_nl;
  wire[22:0] nl_MultLoop_acc_698_nl;
  wire[17:0] MultLoop_acc_697_nl;
  wire[18:0] nl_MultLoop_acc_697_nl;
  wire[23:0] MultLoop_acc_343_nl;
  wire[24:0] nl_MultLoop_acc_343_nl;
  wire[20:0] MultLoop_acc_701_nl;
  wire[22:0] nl_MultLoop_acc_701_nl;
  wire[10:0] MultLoop_acc_1167_nl;
  wire[11:0] nl_MultLoop_acc_1167_nl;
  wire[18:0] MultLoop_acc_1168_nl;
  wire[19:0] nl_MultLoop_acc_1168_nl;
  wire[17:0] MultLoop_acc_711_nl;
  wire[20:0] nl_MultLoop_acc_711_nl;
  wire[20:0] MultLoop_acc_344_nl;
  wire[21:0] nl_MultLoop_acc_344_nl;
  wire[17:0] MultLoop_acc_691_nl;
  wire[18:0] nl_MultLoop_acc_691_nl;
  wire[11:0] MultLoop_acc_1169_nl;
  wire[12:0] nl_MultLoop_acc_1169_nl;
  wire[24:0] MultLoop_acc_188_nl;
  wire[25:0] nl_MultLoop_acc_188_nl;
  wire[20:0] MultLoop_acc_1351_nl;
  wire[21:0] nl_MultLoop_acc_1351_nl;
  wire[14:0] MultLoop_acc_704_nl;
  wire[15:0] nl_MultLoop_acc_704_nl;
  wire[17:0] MultLoop_acc_185_nl;
  wire[18:0] nl_MultLoop_acc_185_nl;
  wire[23:0] MultLoop_acc_184_nl;
  wire[25:0] nl_MultLoop_acc_184_nl;
  wire[17:0] MultLoop_acc_742_nl;
  wire[19:0] nl_MultLoop_acc_742_nl;
  wire[24:0] MultLoop_acc_179_nl;
  wire[26:0] nl_MultLoop_acc_179_nl;
  wire[16:0] MultLoop_152_MultLoop_acc_3_nl;
  wire[17:0] nl_MultLoop_152_MultLoop_acc_3_nl;
  wire[13:0] MultLoop_acc_732_nl;
  wire[14:0] nl_MultLoop_acc_732_nl;
  wire[17:0] MultLoop_acc_1163_nl;
  wire[18:0] nl_MultLoop_acc_1163_nl;
  wire[21:0] MultLoop_acc_730_nl;
  wire[22:0] nl_MultLoop_acc_730_nl;
  wire[12:0] MultLoop_acc_1162_nl;
  wire[13:0] nl_MultLoop_acc_1162_nl;
  wire[18:0] MultLoop_acc_1349_nl;
  wire[19:0] nl_MultLoop_acc_1349_nl;
  wire[18:0] MultLoop_acc_1164_nl;
  wire[19:0] nl_MultLoop_acc_1164_nl;
  wire[23:0] MultLoop_acc_735_nl;
  wire[24:0] nl_MultLoop_acc_735_nl;
  wire[21:0] MultLoop_acc_734_nl;
  wire[22:0] nl_MultLoop_acc_734_nl;
  wire[22:0] MultLoop_acc_340_nl;
  wire[23:0] nl_MultLoop_acc_340_nl;
  wire[17:0] MultLoop_acc_1155_nl;
  wire[18:0] nl_MultLoop_acc_1155_nl;
  wire[24:0] MultLoop_acc_719_nl;
  wire[25:0] nl_MultLoop_acc_719_nl;
  wire[21:0] MultLoop_acc_718_nl;
  wire[23:0] nl_MultLoop_acc_718_nl;
  wire[17:0] MultLoop_acc_1153_nl;
  wire[18:0] nl_MultLoop_acc_1153_nl;
  wire[18:0] MultLoop_acc_1386_nl;
  wire[19:0] nl_MultLoop_acc_1386_nl;
  wire[17:0] MultLoop_acc_1157_nl;
  wire[18:0] nl_MultLoop_acc_1157_nl;
  wire[24:0] MultLoop_acc_722_nl;
  wire[26:0] nl_MultLoop_acc_722_nl;
  wire[17:0] MultLoop_acc_1160_nl;
  wire[18:0] nl_MultLoop_acc_1160_nl;
  wire[18:0] MultLoop_acc_1159_nl;
  wire[19:0] nl_MultLoop_acc_1159_nl;
  wire[22:0] MultLoop_acc_725_nl;
  wire[23:0] nl_MultLoop_acc_725_nl;
  wire[19:0] MultLoop_acc_724_nl;
  wire[20:0] nl_MultLoop_acc_724_nl;
  wire[18:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_4_nl;
  wire[19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_4_nl;
  wire[18:0] MultLoop_acc_594_nl;
  wire[19:0] nl_MultLoop_acc_594_nl;
  wire[17:0] Result_acc_71_nl;
  wire[18:0] nl_Result_acc_71_nl;
  wire[19:0] MultLoop_acc_19_nl;
  wire[20:0] nl_MultLoop_acc_19_nl;
  wire[18:0] MultLoop_acc_395_nl;
  wire[19:0] nl_MultLoop_acc_395_nl;
  wire[14:0] MultLoop_acc_1147_nl;
  wire[15:0] nl_MultLoop_acc_1147_nl;
  wire[22:0] MultLoop_acc_213_nl;
  wire[23:0] nl_MultLoop_acc_213_nl;
  wire[17:0] Result_acc_46_nl;
  wire[18:0] nl_Result_acc_46_nl;
  wire[21:0] MultLoop_acc_123_nl;
  wire[22:0] nl_MultLoop_acc_123_nl;
  wire[20:0] MultLoop_acc_865_nl;
  wire[21:0] nl_MultLoop_acc_865_nl;
  wire[20:0] Result_acc_41_nl;
  wire[21:0] nl_Result_acc_41_nl;
  wire[18:0] Result_acc_138_nl;
  wire[19:0] nl_Result_acc_138_nl;
  wire[13:0] Result_acc_218_nl;
  wire[14:0] nl_Result_acc_218_nl;
  wire[23:0] MultLoop_acc_302_nl;
  wire[24:0] nl_MultLoop_acc_302_nl;
  wire[17:0] MultLoop_acc_397_nl;
  wire[18:0] nl_MultLoop_acc_397_nl;
  wire[22:0] MultLoop_acc_45_nl;
  wire[23:0] nl_MultLoop_acc_45_nl;
  wire[20:0] MultLoop_acc_1049_nl;
  wire[21:0] nl_MultLoop_acc_1049_nl;
  wire[20:0] MultLoop_acc_808_nl;
  wire[21:0] nl_MultLoop_acc_808_nl;
  wire[17:0] MultLoop_acc_56_nl;
  wire[18:0] nl_MultLoop_acc_56_nl;
  wire[17:0] MultLoop_acc_74_nl;
  wire[18:0] nl_MultLoop_acc_74_nl;
  wire[20:0] MultLoop_acc_596_nl;
  wire[21:0] nl_MultLoop_acc_596_nl;
  wire[19:0] MultLoop_acc_714_nl;
  wire[20:0] nl_MultLoop_acc_714_nl;
  wire[20:0] MultLoop_acc_279_nl;
  wire[21:0] nl_MultLoop_acc_279_nl;
  wire[18:0] MultLoop_acc_916_nl;
  wire[19:0] nl_MultLoop_acc_916_nl;
  wire[10:0] MultLoop_acc_1265_nl;
  wire[11:0] nl_MultLoop_acc_1265_nl;
  wire[19:0] MultLoop_acc_694_nl;
  wire[21:0] nl_MultLoop_acc_694_nl;
  wire[18:0] MultLoop_acc_1374_nl;
  wire[19:0] nl_MultLoop_acc_1374_nl;
  wire[10:0] MultLoop_acc_1177_nl;
  wire[11:0] nl_MultLoop_acc_1177_nl;
  wire[22:0] MultLoop_acc_237_nl;
  wire[23:0] nl_MultLoop_acc_237_nl;
  wire[19:0] MultLoop_acc_1354_nl;
  wire[20:0] nl_MultLoop_acc_1354_nl;
  wire[19:0] MultLoop_acc_114_nl;
  wire[20:0] nl_MultLoop_acc_114_nl;
  wire[18:0] MultLoop_acc_404_nl;
  wire[19:0] nl_MultLoop_acc_404_nl;
  wire[17:0] MultLoop_acc_398_nl;
  wire[18:0] nl_MultLoop_acc_398_nl;
  wire[19:0] MultLoop_acc_108_nl;
  wire[20:0] nl_MultLoop_acc_108_nl;
  wire[18:0] MultLoop_acc_402_nl;
  wire[19:0] nl_MultLoop_acc_402_nl;
  wire[13:0] MultLoop_acc_1149_nl;
  wire[14:0] nl_MultLoop_acc_1149_nl;
  wire[23:0] MultLoop_acc_100_nl;
  wire[24:0] nl_MultLoop_acc_100_nl;
  wire[22:0] MultLoop_acc_400_nl;
  wire[23:0] nl_MultLoop_acc_400_nl;
  wire[23:0] MultLoop_acc_554_nl;
  wire[24:0] nl_MultLoop_acc_554_nl;
  wire[22:0] MultLoop_acc_901_nl;
  wire[23:0] nl_MultLoop_acc_901_nl;
  wire[19:0] MultLoop_acc_900_nl;
  wire[20:0] nl_MultLoop_acc_900_nl;
  wire[17:0] MultLoop_acc_899_nl;
  wire[18:0] nl_MultLoop_acc_899_nl;
  wire[9:0] MultLoop_acc_1247_nl;
  wire[10:0] nl_MultLoop_acc_1247_nl;
  wire[18:0] MultLoop_acc_751_nl;
  wire[19:0] nl_MultLoop_acc_751_nl;
  wire[18:0] MultLoop_acc_620_nl;
  wire[19:0] nl_MultLoop_acc_620_nl;
  wire[20:0] MultLoop_acc_130_nl;
  wire[21:0] nl_MultLoop_acc_130_nl;
  wire[16:0] MultLoop_acc_1229_nl;
  wire[17:0] nl_MultLoop_acc_1229_nl;
  wire[18:0] MultLoop_acc_731_nl;
  wire[19:0] nl_MultLoop_acc_731_nl;
  wire[22:0] MultLoop_acc_660_nl;
  wire[23:0] nl_MultLoop_acc_660_nl;
  wire[20:0] MultLoop_acc_206_nl;
  wire[21:0] nl_MultLoop_acc_206_nl;
  wire[17:0] MultLoop_acc_409_nl;
  wire[18:0] nl_MultLoop_acc_409_nl;
  wire[18:0] MultLoop_acc_1198_nl;
  wire[19:0] nl_MultLoop_acc_1198_nl;
  wire[19:0] MultLoop_acc_793_nl;
  wire[20:0] nl_MultLoop_acc_793_nl;
  wire[24:0] MultLoop_acc_159_nl;
  wire[25:0] nl_MultLoop_acc_159_nl;
  wire[23:0] MultLoop_acc_407_nl;
  wire[24:0] nl_MultLoop_acc_407_nl;
  wire[17:0] MultLoop_acc_170_nl;
  wire[18:0] nl_MultLoop_acc_170_nl;
  wire[20:0] MultLoop_acc_1395_nl;
  wire[22:0] nl_MultLoop_acc_1395_nl;
  wire[21:0] MultLoop_acc_1397_nl;
  wire[22:0] nl_MultLoop_acc_1397_nl;
  wire[20:0] MultLoop_acc_1399_nl;
  wire[21:0] nl_MultLoop_acc_1399_nl;
  wire[20:0] MultLoop_acc_1401_nl;
  wire[22:0] nl_MultLoop_acc_1401_nl;
  wire[20:0] MultLoop_acc_1403_nl;
  wire[21:0] nl_MultLoop_acc_1403_nl;
  wire[18:0] MultLoop_acc_1348_nl;
  wire[19:0] nl_MultLoop_acc_1348_nl;
  wire[18:0] MultLoop_acc_1350_nl;
  wire[19:0] nl_MultLoop_acc_1350_nl;
  wire[22:0] MultLoop_acc_353_nl;
  wire[23:0] nl_MultLoop_acc_353_nl;
  wire[19:0] MultLoop_acc_411_nl;
  wire[20:0] nl_MultLoop_acc_411_nl;
  wire[22:0] MultLoop_acc_1390_nl;
  wire[23:0] nl_MultLoop_acc_1390_nl;
  wire[20:0] MultLoop_acc_1359_nl;
  wire[21:0] nl_MultLoop_acc_1359_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [575:0] nl_res_rsci_d;
  assign nl_res_rsci_d = {res_rsci_d_575_558 , res_rsci_d_557_540 , res_rsci_d_539_522
      , res_rsci_d_521_504 , res_rsci_d_503_486 , res_rsci_d_485_468 , res_rsci_d_467_450
      , res_rsci_d_449_432 , res_rsci_d_431_414 , res_rsci_d_413_396 , res_rsci_d_395_378
      , res_rsci_d_377_360 , res_rsci_d_359_342 , res_rsci_d_341_324 , res_rsci_d_323_306
      , res_rsci_d_305_288 , res_rsci_d_287_270 , res_rsci_d_269_252 , res_rsci_d_251_234
      , res_rsci_d_233_216 , res_rsci_d_215_198 , res_rsci_d_197_180 , res_rsci_d_179_162
      , res_rsci_d_161_144 , res_rsci_d_143_126 , res_rsci_d_125_108 , res_rsci_d_107_90
      , res_rsci_d_89_72 , res_rsci_d_71_54 , res_rsci_d_53_36 , res_rsci_d_35_18
      , res_rsci_d_17_0};
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd180)) data_rsci (
      .dat(data_rsc_dat),
      .idat(data_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd2),
  .width(32'sd576)) res_rsci (
      .d(nl_res_rsci_d[575:0]),
      .z(res_rsc_z)
    );
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_4_nl = conv_s2s_18_19(data_rsci_idat[17:0])
      + conv_s2s_16_19(data_rsci_idat[17:2]);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_4_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_4_nl[18:0];
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_4_itm_18_2_1 =
      readslicef_19_17_2((nnet_product_input_t_config2_weight_t_config2_accum_t_acc_4_nl));
  assign nl_Result_acc_175_cse = conv_s2s_18_19(data_rsci_idat[143:126]) + conv_s2s_16_19(data_rsci_idat[143:128]);
  assign Result_acc_175_cse = nl_Result_acc_175_cse[18:0];
  assign nl_MultLoop_acc_594_nl = conv_s2s_18_19(data_rsci_idat[17:0]) + conv_s2s_13_19(data_rsci_idat[17:5]);
  assign MultLoop_acc_594_nl = nl_MultLoop_acc_594_nl[18:0];
  assign MultLoop_acc_594_itm_18_2_1 = readslicef_19_17_2((MultLoop_acc_594_nl));
  assign nl_MultLoop_acc_759_sdt_1 = ({(data_rsci_idat[35:18]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[35:18]));
  assign MultLoop_acc_759_sdt_1 = nl_MultLoop_acc_759_sdt_1[20:0];
  assign nl_Result_acc_71_nl = conv_s2u_16_18(data_rsci_idat[53:38]) - (data_rsci_idat[53:36]);
  assign Result_acc_71_nl = nl_Result_acc_71_nl[17:0];
  assign Result_acc_71_itm_17_7 = readslicef_18_11_7((Result_acc_71_nl));
  assign nl_MultLoop_acc_1254_cse_1 = conv_s2u_11_12(data_rsci_idat[17:7]) + 12'b000000000001;
  assign MultLoop_acc_1254_cse_1 = nl_MultLoop_acc_1254_cse_1[11:0];
  assign nl_MultLoop_acc_1213_cse_1 = conv_s2u_8_9(data_rsci_idat[71:64]) + 9'b000000001;
  assign MultLoop_acc_1213_cse_1 = nl_MultLoop_acc_1213_cse_1[8:0];
  assign nl_MultLoop_acc_1147_nl = conv_s2s_14_15(data_rsci_idat[125:112]) + 15'b000000000000001;
  assign MultLoop_acc_1147_nl = nl_MultLoop_acc_1147_nl[14:0];
  assign nl_MultLoop_acc_395_nl = conv_s2s_18_19(data_rsci_idat[125:108]) + conv_s2s_17_19({(MultLoop_acc_1147_nl)
      , (data_rsci_idat[111:110])});
  assign MultLoop_acc_395_nl = nl_MultLoop_acc_395_nl[18:0];
  assign nl_MultLoop_acc_19_nl = conv_s2u_19_20(MultLoop_acc_395_nl) + ({(~ (data_rsci_idat[125:108]))
      , 2'b00});
  assign MultLoop_acc_19_nl = nl_MultLoop_acc_19_nl[19:0];
  assign MultLoop_acc_19_itm_19_3 = readslicef_20_17_3((MultLoop_acc_19_nl));
  assign nl_MultLoop_acc_1273_cse_1 = conv_s2u_9_10(data_rsci_idat[179:171]) + 10'b0000000001;
  assign MultLoop_acc_1273_cse_1 = nl_MultLoop_acc_1273_cse_1[9:0];
  assign nl_MultLoop_acc_875_cse_1 = conv_s2s_18_19(data_rsci_idat[35:18]) + conv_s2s_16_19(data_rsci_idat[35:20]);
  assign MultLoop_acc_875_cse_1 = nl_MultLoop_acc_875_cse_1[18:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_5_cse_1 = conv_s2s_21_22({(~
      (data_rsci_idat[17:0])) , 3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[17:0]));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_5_cse_1 = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_5_cse_1[21:0];
  assign nl_MultLoop_acc_1148_cse_1 = conv_s2u_11_12(data_rsci_idat[71:61]) + 12'b000000000001;
  assign MultLoop_acc_1148_cse_1 = nl_MultLoop_acc_1148_cse_1[11:0];
  assign nl_MultLoop_acc_634_cse_1 = (~ (data_rsci_idat[179:162])) + conv_s2s_17_18({MultLoop_MultLoop_conc_226_16_4
      , (data_rsci_idat[167:164])});
  assign MultLoop_acc_634_cse_1 = nl_MultLoop_acc_634_cse_1[17:0];
  assign nl_MultLoop_acc_213_nl = conv_s2s_18_23(~ (data_rsci_idat[143:126])) + ({(data_rsci_idat[143:126])
      , 5'b00001});
  assign MultLoop_acc_213_nl = nl_MultLoop_acc_213_nl[22:0];
  assign MultLoop_acc_213_itm_22_7 = readslicef_23_16_7((MultLoop_acc_213_nl));
  assign nl_MultLoop_acc_839_cse_1 = conv_s2s_21_22({(~ (data_rsci_idat[35:18]))
      , 3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[35:18]));
  assign MultLoop_acc_839_cse_1 = nl_MultLoop_acc_839_cse_1[21:0];
  assign nl_MultLoop_acc_892_cse_1 = ({(data_rsci_idat[161:144]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[161:144]));
  assign MultLoop_acc_892_cse_1 = nl_MultLoop_acc_892_cse_1[19:0];
  assign nl_Result_acc_46_nl = conv_s2u_14_18(data_rsci_idat[53:40]) - (data_rsci_idat[53:36]);
  assign Result_acc_46_nl = nl_Result_acc_46_nl[17:0];
  assign Result_acc_46_itm_17_4 = readslicef_18_14_4((Result_acc_46_nl));
  assign nl_MultLoop_acc_865_nl = conv_s2s_20_21({(~ (data_rsci_idat[71:54])) , 2'b01})
      + conv_s2s_18_21(~ (data_rsci_idat[71:54]));
  assign MultLoop_acc_865_nl = nl_MultLoop_acc_865_nl[20:0];
  assign nl_MultLoop_acc_123_nl = conv_s2s_21_22(MultLoop_acc_865_nl) + ({(data_rsci_idat[71:54])
      , 4'b0100});
  assign MultLoop_acc_123_nl = nl_MultLoop_acc_123_nl[21:0];
  assign MultLoop_acc_123_itm_21_6 = readslicef_22_16_6((MultLoop_acc_123_nl));
  assign nl_MultLoop_acc_1203_cse_1 = conv_s2u_8_9(data_rsci_idat[53:46]) + 9'b000000001;
  assign MultLoop_acc_1203_cse_1 = nl_MultLoop_acc_1203_cse_1[8:0];
  assign nl_MultLoop_acc_623_cse_1 = ({(data_rsci_idat[143:126]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[143:126]));
  assign MultLoop_acc_623_cse_1 = nl_MultLoop_acc_623_cse_1[20:0];
  assign nl_Result_acc_218_nl = conv_s2s_13_14(data_rsci_idat[179:167]) + 14'b00000000000001;
  assign Result_acc_218_nl = nl_Result_acc_218_nl[13:0];
  assign nl_Result_acc_138_nl = conv_s2s_18_19(data_rsci_idat[179:162]) + conv_s2s_17_19({(Result_acc_218_nl)
      , (data_rsci_idat[166:164])});
  assign Result_acc_138_nl = nl_Result_acc_138_nl[18:0];
  assign nl_Result_acc_41_nl = conv_s2u_19_21(Result_acc_138_nl) + ({(~ (data_rsci_idat[179:162]))
      , 3'b000});
  assign Result_acc_41_nl = nl_Result_acc_41_nl[20:0];
  assign Result_acc_41_itm_20_8 = readslicef_21_13_8((Result_acc_41_nl));
  assign nl_MultLoop_acc_1178_cse_1 = conv_s2u_12_13(data_rsci_idat[53:42]) + 13'b0000000000001;
  assign MultLoop_acc_1178_cse_1 = nl_MultLoop_acc_1178_cse_1[12:0];
  assign nl_MultLoop_acc_565_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[161:144]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[161:144]));
  assign MultLoop_acc_565_cse_1 = nl_MultLoop_acc_565_cse_1[20:0];
  assign nl_MultLoop_acc_777_sdt_1 = ({(data_rsci_idat[179:162]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[179:162]));
  assign MultLoop_acc_777_sdt_1 = nl_MultLoop_acc_777_sdt_1[19:0];
  assign nl_Result_acc_207_cse_1 = conv_s2u_11_12(data_rsci_idat[125:115]) + 12'b000000000001;
  assign Result_acc_207_cse_1 = nl_Result_acc_207_cse_1[11:0];
  assign nl_MultLoop_acc_397_nl = (~ (data_rsci_idat[71:54])) + conv_s2s_17_18({MultLoop_acc_1148_cse_1
      , (data_rsci_idat[60:56])});
  assign MultLoop_acc_397_nl = nl_MultLoop_acc_397_nl[17:0];
  assign nl_MultLoop_acc_302_nl = conv_s2u_18_24(MultLoop_acc_397_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[71:54])) , 5'b00001});
  assign MultLoop_acc_302_nl = nl_MultLoop_acc_302_nl[23:0];
  assign MultLoop_acc_302_itm_23_7 = readslicef_24_17_7((MultLoop_acc_302_nl));
  assign nl_MultLoop_acc_1049_nl = ({(data_rsci_idat[17:0]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_206_18_5
      , (~ (data_rsci_idat[4:0]))});
  assign MultLoop_acc_1049_nl = nl_MultLoop_acc_1049_nl[20:0];
  assign nl_MultLoop_acc_45_nl = conv_s2s_21_23(MultLoop_acc_1049_nl) + ({(~ (data_rsci_idat[17:0]))
      , 5'b00000});
  assign MultLoop_acc_45_nl = nl_MultLoop_acc_45_nl[22:0];
  assign MultLoop_acc_45_itm_22_9 = readslicef_23_14_9((MultLoop_acc_45_nl));
  assign nl_MultLoop_acc_543_cse_1 = (~ (data_rsci_idat[35:18])) + conv_s2s_16_18(data_rsci_idat[35:20]);
  assign MultLoop_acc_543_cse_1 = nl_MultLoop_acc_543_cse_1[17:0];
  assign nl_MultLoop_acc_1017_cse_1 = (~ (data_rsci_idat[89:72])) + conv_s2s_16_18(data_rsci_idat[89:74]);
  assign MultLoop_acc_1017_cse_1 = nl_MultLoop_acc_1017_cse_1[17:0];
  assign nl_MultLoop_acc_405_cse_1 = conv_s2s_18_19(data_rsci_idat[107:90]) + conv_s2s_16_19(data_rsci_idat[107:92]);
  assign MultLoop_acc_405_cse_1 = nl_MultLoop_acc_405_cse_1[18:0];
  assign nl_MultLoop_acc_473_cse_1 = conv_s2s_21_22({(~ (data_rsci_idat[71:54]))
      , 3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[71:54]));
  assign MultLoop_acc_473_cse_1 = nl_MultLoop_acc_473_cse_1[21:0];
  assign nl_MultLoop_acc_763_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[161:144]))
      , 2'b01}) + conv_s2s_19_21({MultLoop_MultLoop_conc_208_18_8 , (~ (data_rsci_idat[151:144]))});
  assign MultLoop_acc_763_cse_1 = nl_MultLoop_acc_763_cse_1[20:0];
  assign nl_Result_acc_202_cse_1 = conv_s2u_9_10(data_rsci_idat[143:135]) + 10'b0000000001;
  assign Result_acc_202_cse_1 = nl_Result_acc_202_cse_1[9:0];
  assign nl_Result_acc_195_cse_1 = (~ (data_rsci_idat[179:162])) + conv_s2s_16_18(data_rsci_idat[179:164]);
  assign Result_acc_195_cse_1 = nl_Result_acc_195_cse_1[17:0];
  assign nl_MultLoop_acc_650_cse_1 = conv_s2s_18_19(data_rsci_idat[125:108]) + conv_s2s_16_19(data_rsci_idat[125:110]);
  assign MultLoop_acc_650_cse_1 = nl_MultLoop_acc_650_cse_1[18:0];
  assign nl_MultLoop_acc_1151_cse_1 = conv_s2u_10_11(data_rsci_idat[17:8]) + 11'b00000000001;
  assign MultLoop_acc_1151_cse_1 = nl_MultLoop_acc_1151_cse_1[10:0];
  assign nl_MultLoop_acc_557_cse_1 = (~ (data_rsci_idat[35:18])) + conv_s2s_15_18(data_rsci_idat[35:21]);
  assign MultLoop_acc_557_cse_1 = nl_MultLoop_acc_557_cse_1[17:0];
  assign nl_MultLoop_acc_808_nl = conv_s2s_20_21({(~ (data_rsci_idat[125:108])) ,
      2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[125:108]));
  assign MultLoop_acc_808_nl = nl_MultLoop_acc_808_nl[20:0];
  assign MultLoop_acc_808_itm_20_2_1 = readslicef_21_19_2((MultLoop_acc_808_nl));
  assign nl_MultLoop_acc_789_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[53:36]))
      , 2'b01}) + conv_s2s_19_21({MultLoop_MultLoop_conc_218_18_8 , (~ (data_rsci_idat[43:36]))});
  assign MultLoop_acc_789_cse_1 = nl_MultLoop_acc_789_cse_1[20:0];
  assign nl_MultLoop_acc_56_nl = conv_s2u_16_18(data_rsci_idat[17:2]) - (data_rsci_idat[17:0]);
  assign MultLoop_acc_56_nl = nl_MultLoop_acc_56_nl[17:0];
  assign MultLoop_acc_56_itm_17_1 = readslicef_18_17_1((MultLoop_acc_56_nl));
  assign nl_MultLoop_acc_412_cse_1 = (~ (data_rsci_idat[17:0])) + conv_s2s_15_18(data_rsci_idat[17:3]);
  assign MultLoop_acc_412_cse_1 = nl_MultLoop_acc_412_cse_1[17:0];
  assign nl_MultLoop_acc_1150_cse_1 = conv_s2u_10_11(data_rsci_idat[89:80]) + 11'b00000000001;
  assign MultLoop_acc_1150_cse_1 = nl_MultLoop_acc_1150_cse_1[10:0];
  assign nl_MultLoop_acc_410_cse_1 = (~ (data_rsci_idat[71:54])) + conv_s2s_14_18(data_rsci_idat[71:58]);
  assign MultLoop_acc_410_cse_1 = nl_MultLoop_acc_410_cse_1[17:0];
  assign nl_MultLoop_acc_74_nl = conv_s2u_15_18(data_rsci_idat[143:129]) - (data_rsci_idat[143:126]);
  assign MultLoop_acc_74_nl = nl_MultLoop_acc_74_nl[17:0];
  assign MultLoop_acc_74_itm_17_1 = readslicef_18_17_1((MultLoop_acc_74_nl));
  assign nl_MultLoop_acc_744_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[17:0])) ,
      2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[17:0]));
  assign MultLoop_acc_744_cse_1 = nl_MultLoop_acc_744_cse_1[20:0];
  assign nl_MultLoop_acc_596_nl = ({(data_rsci_idat[53:36]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[53:36]));
  assign MultLoop_acc_596_nl = nl_MultLoop_acc_596_nl[20:0];
  assign MultLoop_acc_596_itm_20_5 = readslicef_21_16_5((MultLoop_acc_596_nl));
  assign nl_MultLoop_acc_714_nl = ({(data_rsci_idat[161:144]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_208_18_8
      , (~ (data_rsci_idat[151:144]))});
  assign MultLoop_acc_714_nl = nl_MultLoop_acc_714_nl[19:0];
  assign MultLoop_acc_714_itm_19_4 = readslicef_20_16_4((MultLoop_acc_714_nl));
  assign nl_MultLoop_acc_733_cse_1 = ({(data_rsci_idat[53:36]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[53:36]));
  assign MultLoop_acc_733_cse_1 = nl_MultLoop_acc_733_cse_1[19:0];
  assign nl_MultLoop_acc_279_nl = conv_s2u_18_21(MultLoop_acc_412_cse_1) + ({(data_rsci_idat[17:0])
      , 3'b001});
  assign MultLoop_acc_279_nl = nl_MultLoop_acc_279_nl[20:0];
  assign MultLoop_acc_279_itm_20_6 = readslicef_21_15_6((MultLoop_acc_279_nl));
  assign nl_MultLoop_acc_1265_nl = conv_s2s_10_11(data_rsci_idat[143:134]) + 11'b00000000001;
  assign MultLoop_acc_1265_nl = nl_MultLoop_acc_1265_nl[10:0];
  assign nl_MultLoop_acc_916_nl = conv_s2s_18_19(data_rsci_idat[143:126]) + conv_s2s_17_19({(MultLoop_acc_1265_nl)
      , (data_rsci_idat[133:128])});
  assign MultLoop_acc_916_nl = nl_MultLoop_acc_916_nl[18:0];
  assign MultLoop_acc_916_itm_18_3 = readslicef_19_16_3((MultLoop_acc_916_nl));
  assign nl_MultLoop_acc_694_nl = ({(~ (data_rsci_idat[71:54])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[71:54])
      + conv_s2s_16_20(data_rsci_idat[71:56]);
  assign MultLoop_acc_694_nl = nl_MultLoop_acc_694_nl[19:0];
  assign MultLoop_acc_694_itm_19_2_1 = readslicef_20_18_2((MultLoop_acc_694_nl));
  assign nl_MultLoop_acc_805_cse_1 = ({(data_rsci_idat[17:0]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[17:0]));
  assign MultLoop_acc_805_cse_1 = nl_MultLoop_acc_805_cse_1[19:0];
  assign nl_MultLoop_acc_1374_nl = conv_s2u_18_19(data_rsci_idat[161:144]) + conv_s2u_16_19(MultLoop_acc_892_cse_1[19:4]);
  assign MultLoop_acc_1374_nl = nl_MultLoop_acc_1374_nl[18:0];
  assign MultLoop_acc_1374_itm_18_1 = readslicef_19_18_1((MultLoop_acc_1374_nl));
  assign nl_MultLoop_acc_1177_nl = conv_s2s_10_11(data_rsci_idat[107:98]) + 11'b00000000001;
  assign MultLoop_acc_1177_nl = nl_MultLoop_acc_1177_nl[10:0];
  assign nl_MultLoop_acc_753_cse_1 = conv_s2s_18_19(data_rsci_idat[107:90]) + conv_s2s_17_19({(MultLoop_acc_1177_nl)
      , (data_rsci_idat[97:92])});
  assign MultLoop_acc_753_cse_1 = nl_MultLoop_acc_753_cse_1[18:0];
  assign nl_MultLoop_acc_786_cse_1 = ({(data_rsci_idat[89:72]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[89:72]));
  assign MultLoop_acc_786_cse_1 = nl_MultLoop_acc_786_cse_1[19:0];
  assign nl_MultLoop_acc_406_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[143:126]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[143:126]));
  assign MultLoop_acc_406_cse_1 = nl_MultLoop_acc_406_cse_1[20:0];
  assign nl_MultLoop_acc_237_nl = conv_s2s_18_23(~ (data_rsci_idat[17:0])) + ({(data_rsci_idat[17:0])
      , 5'b00001});
  assign MultLoop_acc_237_nl = nl_MultLoop_acc_237_nl[22:0];
  assign MultLoop_acc_237_itm_22_9 = readslicef_23_14_9((MultLoop_acc_237_nl));
  assign nl_MultLoop_acc_812_cse_1 = conv_s2s_18_19(data_rsci_idat[35:18]) + conv_s2s_14_19(data_rsci_idat[35:22]);
  assign MultLoop_acc_812_cse_1 = nl_MultLoop_acc_812_cse_1[18:0];
  assign nl_MultLoop_acc_621_cse_1 = (~ (data_rsci_idat[125:108])) + conv_s2s_15_18(data_rsci_idat[125:111]);
  assign MultLoop_acc_621_cse_1 = nl_MultLoop_acc_621_cse_1[17:0];
  assign nl_MultLoop_acc_1354_nl = ({(data_rsci_idat[89:72]) , 2'b01}) + conv_s2u_19_20(MultLoop_acc_745_cse_1[20:2]);
  assign MultLoop_acc_1354_nl = nl_MultLoop_acc_1354_nl[19:0];
  assign MultLoop_acc_1354_itm_19_3 = readslicef_20_17_3((MultLoop_acc_1354_nl));
  assign nl_MultLoop_acc_404_nl = conv_s2s_18_19(data_rsci_idat[89:72]) + conv_s2s_13_19({MultLoop_acc_1150_cse_1
      , (data_rsci_idat[79:78])});
  assign MultLoop_acc_404_nl = nl_MultLoop_acc_404_nl[18:0];
  assign nl_MultLoop_acc_114_nl = conv_s2u_19_20(MultLoop_acc_404_nl) + ({(~ (data_rsci_idat[89:72]))
      , 2'b00});
  assign MultLoop_acc_114_nl = nl_MultLoop_acc_114_nl[19:0];
  assign MultLoop_acc_114_itm_19_3 = readslicef_20_17_3((MultLoop_acc_114_nl));
  assign nl_MultLoop_acc_398_nl = (~ (data_rsci_idat[17:0])) + conv_s2s_16_18(data_rsci_idat[17:2]);
  assign MultLoop_acc_398_nl = nl_MultLoop_acc_398_nl[17:0];
  assign nl_MultLoop_acc_399_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[17:0])) ,
      2'b01}) + conv_s2s_18_21(MultLoop_acc_398_nl);
  assign MultLoop_acc_399_cse_1 = nl_MultLoop_acc_399_cse_1[20:0];
  assign nl_MultLoop_acc_560_cse_1 = conv_s2s_21_22({(~ (data_rsci_idat[53:36]))
      , 3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[53:36]));
  assign MultLoop_acc_560_cse_1 = nl_MultLoop_acc_560_cse_1[21:0];
  assign nl_MultLoop_acc_702_cse_1 = conv_s2s_18_19(data_rsci_idat[179:162]) + conv_s2s_16_19(data_rsci_idat[179:164]);
  assign MultLoop_acc_702_cse_1 = nl_MultLoop_acc_702_cse_1[18:0];
  assign nl_MultLoop_acc_1149_nl = conv_s2s_13_14(data_rsci_idat[161:149]) + 14'b00000000000001;
  assign MultLoop_acc_1149_nl = nl_MultLoop_acc_1149_nl[13:0];
  assign nl_MultLoop_acc_402_nl = conv_s2s_18_19(data_rsci_idat[161:144]) + conv_s2s_16_19({(MultLoop_acc_1149_nl)
      , (data_rsci_idat[148:147])});
  assign MultLoop_acc_402_nl = nl_MultLoop_acc_402_nl[18:0];
  assign nl_MultLoop_acc_108_nl = conv_s2u_19_20(MultLoop_acc_402_nl) + ({(~ (data_rsci_idat[161:144]))
      , 2'b00});
  assign MultLoop_acc_108_nl = nl_MultLoop_acc_108_nl[19:0];
  assign MultLoop_acc_108_itm_19_6 = readslicef_20_14_6((MultLoop_acc_108_nl));
  assign nl_MultLoop_acc_400_nl = conv_s2s_22_23({(~ (data_rsci_idat[17:0])) , 4'b0100})
      + conv_s2s_21_23(MultLoop_acc_399_cse_1);
  assign MultLoop_acc_400_nl = nl_MultLoop_acc_400_nl[22:0];
  assign nl_MultLoop_acc_100_nl = conv_s2u_23_24(MultLoop_acc_400_nl) + ({(data_rsci_idat[17:0])
      , 6'b010000});
  assign MultLoop_acc_100_nl = nl_MultLoop_acc_100_nl[23:0];
  assign MultLoop_acc_100_itm_23_7 = readslicef_24_17_7((MultLoop_acc_100_nl));
  assign nl_MultLoop_acc_745_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[89:72]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[89:72]));
  assign MultLoop_acc_745_cse_1 = nl_MultLoop_acc_745_cse_1[20:0];
  assign nl_MultLoop_acc_1239_cse_1 = conv_s2u_13_14(data_rsci_idat[17:5]) + 14'b00000000000001;
  assign MultLoop_acc_1239_cse_1 = nl_MultLoop_acc_1239_cse_1[13:0];
  assign nl_MultLoop_acc_554_nl = conv_s2s_23_24({(~ (data_rsci_idat[107:90])) ,
      5'b00001}) + conv_s2s_18_24(~ (data_rsci_idat[107:90]));
  assign MultLoop_acc_554_nl = nl_MultLoop_acc_554_nl[23:0];
  assign MultLoop_acc_554_itm_23_5_1 = readslicef_24_19_5((MultLoop_acc_554_nl));
  assign nl_MultLoop_acc_1247_nl = conv_s2s_9_10(data_rsci_idat[53:45]) + 10'b0000000001;
  assign MultLoop_acc_1247_nl = nl_MultLoop_acc_1247_nl[9:0];
  assign nl_MultLoop_acc_899_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_16_18({(MultLoop_acc_1247_nl)
      , (data_rsci_idat[44:39])});
  assign MultLoop_acc_899_nl = nl_MultLoop_acc_899_nl[17:0];
  assign nl_MultLoop_acc_900_nl = ({(data_rsci_idat[53:36]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_899_nl);
  assign MultLoop_acc_900_nl = nl_MultLoop_acc_900_nl[19:0];
  assign nl_MultLoop_acc_901_nl = conv_s2u_22_23({(data_rsci_idat[53:36]) , 4'b0000})
      + conv_s2u_20_23(MultLoop_acc_900_nl);
  assign MultLoop_acc_901_nl = nl_MultLoop_acc_901_nl[22:0];
  assign MultLoop_acc_901_itm_22_5 = readslicef_23_18_5((MultLoop_acc_901_nl));
  assign nl_MultLoop_acc_847_cse_1 = (~ (data_rsci_idat[125:108])) + conv_s2s_16_18(data_rsci_idat[125:110]);
  assign MultLoop_acc_847_cse_1 = nl_MultLoop_acc_847_cse_1[17:0];
  assign nl_MultLoop_acc_751_nl = conv_s2s_18_19(data_rsci_idat[125:108]) + conv_s2s_14_19(data_rsci_idat[125:112]);
  assign MultLoop_acc_751_nl = nl_MultLoop_acc_751_nl[18:0];
  assign MultLoop_acc_751_itm_18_2 = readslicef_19_17_2((MultLoop_acc_751_nl));
  assign nl_MultLoop_acc_578_cse_1 = conv_s2s_21_22({(~ (data_rsci_idat[89:72]))
      , 3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[89:72]));
  assign MultLoop_acc_578_cse_1 = nl_MultLoop_acc_578_cse_1[21:0];
  assign nl_MultLoop_acc_620_nl = conv_s2s_18_19(data_rsci_idat[107:90]) + conv_s2s_14_19(data_rsci_idat[107:94]);
  assign MultLoop_acc_620_nl = nl_MultLoop_acc_620_nl[18:0];
  assign MultLoop_acc_620_itm_18_3 = readslicef_19_16_3((MultLoop_acc_620_nl));
  assign nl_MultLoop_acc_642_cse_1 = (~ (data_rsci_idat[53:36])) + conv_s2s_14_18({MultLoop_acc_1203_cse_1
      , (data_rsci_idat[45:41])});
  assign MultLoop_acc_642_cse_1 = nl_MultLoop_acc_642_cse_1[17:0];
  assign nl_MultLoop_acc_1229_nl =  -conv_s2s_16_17(data_rsci_idat[17:2]);
  assign MultLoop_acc_1229_nl = nl_MultLoop_acc_1229_nl[16:0];
  assign nl_MultLoop_acc_130_nl = conv_s2s_19_21({(MultLoop_acc_1229_nl) , (~ (data_rsci_idat[1:0]))})
      + conv_s2s_20_21({(~ (data_rsci_idat[17:0])) , 2'b01});
  assign MultLoop_acc_130_nl = nl_MultLoop_acc_130_nl[20:0];
  assign MultLoop_acc_130_itm_20_10 = readslicef_21_11_10((MultLoop_acc_130_nl));
  assign nl_MultLoop_acc_731_nl = conv_s2s_18_19(data_rsci_idat[17:0]) + conv_s2s_15_19(data_rsci_idat[17:3]);
  assign MultLoop_acc_731_nl = nl_MultLoop_acc_731_nl[18:0];
  assign MultLoop_acc_731_itm_18_4 = readslicef_19_15_4((MultLoop_acc_731_nl));
  assign nl_MultLoop_acc_660_nl = conv_s2s_22_23({(~ (data_rsci_idat[89:72])) , 4'b0001})
      + conv_s2s_18_23(~ (data_rsci_idat[89:72]));
  assign MultLoop_acc_660_nl = nl_MultLoop_acc_660_nl[22:0];
  assign MultLoop_acc_660_itm_22_4_1 = readslicef_23_19_4((MultLoop_acc_660_nl));
  assign nl_MultLoop_acc_409_nl = (~ (data_rsci_idat[17:0])) + conv_s2s_13_18({MultLoop_acc_1151_cse_1
      , (data_rsci_idat[7:6])});
  assign MultLoop_acc_409_nl = nl_MultLoop_acc_409_nl[17:0];
  assign nl_MultLoop_acc_206_nl = conv_s2u_18_21(MultLoop_acc_409_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[17:0])) , 2'b01});
  assign MultLoop_acc_206_nl = nl_MultLoop_acc_206_nl[20:0];
  assign MultLoop_acc_206_itm_20_4 = readslicef_21_17_4((MultLoop_acc_206_nl));
  assign nl_MultLoop_acc_793_nl = ({(data_rsci_idat[161:144]) , 2'b01}) + conv_s2s_19_20({Result_Result_conc_52_18_10
      , (~ (data_rsci_idat[153:144]))});
  assign MultLoop_acc_793_nl = nl_MultLoop_acc_793_nl[19:0];
  assign nl_MultLoop_acc_1198_nl = conv_s2u_18_19(data_rsci_idat[161:144]) + conv_s2u_13_19(readslicef_20_13_7((MultLoop_acc_793_nl)));
  assign MultLoop_acc_1198_nl = nl_MultLoop_acc_1198_nl[18:0];
  assign MultLoop_acc_1198_itm_18_2 = readslicef_19_17_2((MultLoop_acc_1198_nl));
  assign nl_MultLoop_acc_407_nl = conv_s2s_23_24({(~ (data_rsci_idat[143:126])) ,
      5'b00100}) + conv_s2s_21_24(MultLoop_acc_406_cse_1);
  assign MultLoop_acc_407_nl = nl_MultLoop_acc_407_nl[23:0];
  assign nl_MultLoop_acc_159_nl = conv_s2s_24_25(MultLoop_acc_407_nl) + ({(data_rsci_idat[143:126])
      , 7'b0100000});
  assign MultLoop_acc_159_nl = nl_MultLoop_acc_159_nl[24:0];
  assign MultLoop_acc_159_itm_24_9 = readslicef_25_16_9((MultLoop_acc_159_nl));
  assign nl_MultLoop_acc_170_nl = conv_s2u_16_18(data_rsci_idat[143:128]) - (data_rsci_idat[143:126]);
  assign MultLoop_acc_170_nl = nl_MultLoop_acc_170_nl[17:0];
  assign MultLoop_acc_170_itm_17_8 = readslicef_18_10_8((MultLoop_acc_170_nl));
  assign nl_Result_Result_conc_48_18_9 =  -conv_s2s_9_10(data_rsci_idat[143:135]);
  assign Result_Result_conc_48_18_9 = nl_Result_Result_conc_48_18_9[9:0];
  assign nl_MultLoop_MultLoop_conc_202_18_7 =  -conv_s2s_11_12(data_rsci_idat[71:61]);
  assign MultLoop_MultLoop_conc_202_18_7 = nl_MultLoop_MultLoop_conc_202_18_7[11:0];
  assign nl_MultLoop_acc_1395_nl = ({(~ (data_rsci_idat[53:36])) , 3'b000}) + conv_s2s_18_21(data_rsci_idat[53:36])
      + conv_s2s_15_21(data_rsci_idat[53:39]);
  assign MultLoop_acc_1395_nl = nl_MultLoop_acc_1395_nl[20:0];
  assign MultLoop_acc_1395_itm_20_3_1 = readslicef_21_18_3((MultLoop_acc_1395_nl));
  assign nl_Result_Result_conc_50_13_2 = conv_s2s_11_12(data_rsci_idat[53:43]) +
      12'b000000000001;
  assign Result_Result_conc_50_13_2 = nl_Result_Result_conc_50_13_2[11:0];
  assign nl_MultLoop_MultLoop_conc_204_18_9 =  -conv_s2s_9_10(data_rsci_idat[89:81]);
  assign MultLoop_MultLoop_conc_204_18_9 = nl_MultLoop_MultLoop_conc_204_18_9[9:0];
  assign nl_Result_Result_conc_52_18_10 =  -conv_s2s_8_9(data_rsci_idat[161:154]);
  assign Result_Result_conc_52_18_10 = nl_Result_Result_conc_52_18_10[8:0];
  assign nl_Result_Result_conc_54_18_8 =  -conv_s2s_10_11(data_rsci_idat[89:80]);
  assign Result_Result_conc_54_18_8 = nl_Result_Result_conc_54_18_8[10:0];
  assign nl_MultLoop_MultLoop_conc_206_18_5 =  -conv_s2s_13_14(data_rsci_idat[17:5]);
  assign MultLoop_MultLoop_conc_206_18_5 = nl_MultLoop_MultLoop_conc_206_18_5[13:0];
  assign nl_MultLoop_acc_1397_nl = conv_s2s_21_22({(~ (data_rsci_idat[71:54])) ,
      3'b001}) + conv_s2s_19_22({MultLoop_MultLoop_conc_202_18_7 , (~ (data_rsci_idat[60:54]))});
  assign MultLoop_acc_1397_nl = nl_MultLoop_acc_1397_nl[21:0];
  assign MultLoop_acc_1397_itm_21_3_1 = readslicef_22_19_3((MultLoop_acc_1397_nl));
  assign nl_MultLoop_MultLoop_conc_208_18_8 =  -conv_s2s_10_11(data_rsci_idat[161:152]);
  assign MultLoop_MultLoop_conc_208_18_8 = nl_MultLoop_MultLoop_conc_208_18_8[10:0];
  assign nl_Result_Result_conc_56_18_6 =  -conv_s2s_12_13(data_rsci_idat[89:78]);
  assign Result_Result_conc_56_18_6 = nl_Result_Result_conc_56_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_210_18_8 =  -conv_s2s_10_11(data_rsci_idat[35:26]);
  assign MultLoop_MultLoop_conc_210_18_8 = nl_MultLoop_MultLoop_conc_210_18_8[10:0];
  assign nl_Result_Result_conc_58_18_9 =  -conv_s2s_9_10(data_rsci_idat[107:99]);
  assign Result_Result_conc_58_18_9 = nl_Result_Result_conc_58_18_9[9:0];
  assign nl_MultLoop_MultLoop_conc_212_18_6 =  -conv_s2s_12_13(data_rsci_idat[161:150]);
  assign MultLoop_MultLoop_conc_212_18_6 = nl_MultLoop_MultLoop_conc_212_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_214_18_10 =  -conv_s2s_8_9(data_rsci_idat[53:46]);
  assign MultLoop_MultLoop_conc_214_18_10 = nl_MultLoop_MultLoop_conc_214_18_10[8:0];
  assign nl_Result_Result_conc_60_18_7 =  -conv_s2s_11_12(data_rsci_idat[107:97]);
  assign Result_Result_conc_60_18_7 = nl_Result_Result_conc_60_18_7[11:0];
  assign nl_MultLoop_acc_1399_nl = ({(data_rsci_idat[89:72]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_204_18_9
      , (~ (data_rsci_idat[80:72]))});
  assign MultLoop_acc_1399_nl = nl_MultLoop_acc_1399_nl[20:0];
  assign MultLoop_acc_1399_itm_20_5 = readslicef_21_16_5((MultLoop_acc_1399_nl));
  assign nl_MultLoop_MultLoop_conc_216_18_8 =  -conv_s2s_10_11(data_rsci_idat[179:170]);
  assign MultLoop_MultLoop_conc_216_18_8 = nl_MultLoop_MultLoop_conc_216_18_8[10:0];
  assign nl_Result_Result_conc_62_18_6 =  -conv_s2s_12_13(data_rsci_idat[107:96]);
  assign Result_Result_conc_62_18_6 = nl_Result_Result_conc_62_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_218_18_8 =  -conv_s2s_10_11(data_rsci_idat[53:44]);
  assign MultLoop_MultLoop_conc_218_18_8 = nl_MultLoop_MultLoop_conc_218_18_8[10:0];
  assign nl_MultLoop_acc_1401_nl = conv_s2s_20_21({(data_rsci_idat[161:144]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[161:144]) + conv_s2s_16_21(data_rsci_idat[161:146]);
  assign MultLoop_acc_1401_nl = nl_MultLoop_acc_1401_nl[20:0];
  assign MultLoop_acc_1401_itm_20_5 = readslicef_21_16_5((MultLoop_acc_1401_nl));
  assign nl_MultLoop_MultLoop_conc_222_18_9 =  -conv_s2s_9_10(data_rsci_idat[125:117]);
  assign MultLoop_MultLoop_conc_222_18_9 = nl_MultLoop_MultLoop_conc_222_18_9[9:0];
  assign nl_MultLoop_MultLoop_conc_224_16_6 = conv_s2s_10_11(data_rsci_idat[179:170])
      + 11'b00000000001;
  assign MultLoop_MultLoop_conc_224_16_6 = nl_MultLoop_MultLoop_conc_224_16_6[10:0];
  assign nl_MultLoop_acc_1403_nl = conv_s2s_20_21({(~ (data_rsci_idat[35:18])) ,
      2'b01}) + conv_s2s_18_21(MultLoop_acc_543_cse_1);
  assign MultLoop_acc_1403_nl = nl_MultLoop_acc_1403_nl[20:0];
  assign MultLoop_acc_1403_itm_20_2_1 = readslicef_21_19_2((MultLoop_acc_1403_nl));
  assign nl_MultLoop_MultLoop_conc_226_16_4 = conv_s2s_12_13(data_rsci_idat[179:168])
      + 13'b0000000000001;
  assign MultLoop_MultLoop_conc_226_16_4 = nl_MultLoop_MultLoop_conc_226_16_4[12:0];
  assign nl_MultLoop_MultLoop_conc_228_18_9 =  -conv_s2s_9_10(data_rsci_idat[71:63]);
  assign MultLoop_MultLoop_conc_228_18_9 = nl_MultLoop_MultLoop_conc_228_18_9[9:0];
  assign nl_Result_Result_conc_64_18_8 =  -conv_s2s_10_11(data_rsci_idat[71:62]);
  assign Result_Result_conc_64_18_8 = nl_Result_Result_conc_64_18_8[10:0];
  assign nl_MultLoop_acc_1348_nl = conv_s2u_16_19(MultLoop_acc_405_cse_1[18:3]) +
      conv_s2u_18_19(data_rsci_idat[107:90]);
  assign MultLoop_acc_1348_nl = nl_MultLoop_acc_1348_nl[18:0];
  assign MultLoop_acc_1348_itm_18_3 = readslicef_19_16_3((MultLoop_acc_1348_nl));
  assign nl_MultLoop_acc_1350_nl = conv_s2u_18_19(data_rsci_idat[179:162]) + conv_s2u_17_19(MultLoop_acc_702_cse_1[18:2]);
  assign MultLoop_acc_1350_nl = nl_MultLoop_acc_1350_nl[18:0];
  assign MultLoop_acc_1350_itm_18_5 = readslicef_19_14_5((MultLoop_acc_1350_nl));
  assign nl_MultLoop_acc_411_nl = ({(data_rsci_idat[71:54]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_410_cse_1);
  assign MultLoop_acc_411_nl = nl_MultLoop_acc_411_nl[19:0];
  assign nl_MultLoop_acc_353_nl = conv_s2u_20_23(MultLoop_acc_411_nl) + conv_s2u_22_23({(data_rsci_idat[71:54])
      , 4'b0000});
  assign MultLoop_acc_353_nl = nl_MultLoop_acc_353_nl[22:0];
  assign MultLoop_acc_353_itm_22_6 = readslicef_23_17_6((MultLoop_acc_353_nl));
  assign nl_MultLoop_acc_1390_nl = conv_s2u_22_23({(~ (data_rsci_idat[161:144]))
      , 4'b0001}) + conv_s2u_19_23(MultLoop_acc_565_cse_1[20:2]);
  assign MultLoop_acc_1390_nl = nl_MultLoop_acc_1390_nl[22:0];
  assign MultLoop_acc_1390_itm_22_4_1 = readslicef_23_19_4((MultLoop_acc_1390_nl));
  assign nl_MultLoop_asn_361 = (~ (data_rsci_idat[179:162])) + conv_s2s_17_18(MultLoop_acc_702_cse_1[18:2]);
  assign MultLoop_asn_361 = nl_MultLoop_asn_361[17:0];
  assign nl_MultLoop_acc_1359_nl = conv_s2u_20_21({(~ (data_rsci_idat[125:108]))
      , 2'b01}) + conv_s2u_19_21(MultLoop_acc_808_itm_20_2_1);
  assign MultLoop_acc_1359_nl = nl_MultLoop_acc_1359_nl[20:0];
  assign MultLoop_acc_1359_itm_20_2_1 = readslicef_21_19_2((MultLoop_acc_1359_nl));
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      res_rsci_d_575_558 <= 18'b000000000000000000;
      res_rsci_d_17_0 <= 18'b000000000000000000;
      res_rsci_d_557_540 <= 18'b000000000000000000;
      res_rsci_d_35_18 <= 18'b000000000000000000;
      res_rsci_d_539_522 <= 18'b000000000000000000;
      res_rsci_d_53_36 <= 18'b000000000000000000;
      res_rsci_d_521_504 <= 18'b000000000000000000;
      res_rsci_d_71_54 <= 18'b000000000000000000;
      res_rsci_d_503_486 <= 18'b000000000000000000;
      res_rsci_d_89_72 <= 18'b000000000000000000;
      res_rsci_d_485_468 <= 18'b000000000000000000;
      res_rsci_d_107_90 <= 18'b000000000000000000;
      res_rsci_d_467_450 <= 18'b000000000000000000;
      res_rsci_d_125_108 <= 18'b000000000000000000;
      res_rsci_d_449_432 <= 18'b000000000000000000;
      res_rsci_d_143_126 <= 18'b000000000000000000;
      res_rsci_d_431_414 <= 18'b000000000000000000;
      res_rsci_d_161_144 <= 18'b000000000000000000;
      res_rsci_d_413_396 <= 18'b000000000000000000;
      res_rsci_d_179_162 <= 18'b000000000000000000;
      res_rsci_d_395_378 <= 18'b000000000000000000;
      res_rsci_d_197_180 <= 18'b000000000000000000;
      res_rsci_d_377_360 <= 18'b000000000000000000;
      res_rsci_d_215_198 <= 18'b000000000000000000;
      res_rsci_d_359_342 <= 18'b000000000000000000;
      res_rsci_d_233_216 <= 18'b000000000000000000;
      res_rsci_d_341_324 <= 18'b000000000000000000;
      res_rsci_d_251_234 <= 18'b000000000000000000;
      res_rsci_d_323_306 <= 18'b000000000000000000;
      res_rsci_d_269_252 <= 18'b000000000000000000;
      res_rsci_d_305_288 <= 18'b000000000000000000;
      res_rsci_d_287_270 <= 18'b000000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      res_rsci_d_575_558 <= nl_res_rsci_d_575_558[17:0];
      res_rsci_d_17_0 <= nl_res_rsci_d_17_0[17:0];
      res_rsci_d_557_540 <= nl_res_rsci_d_557_540[17:0];
      res_rsci_d_35_18 <= nl_res_rsci_d_35_18[17:0];
      res_rsci_d_539_522 <= nl_res_rsci_d_539_522[17:0];
      res_rsci_d_53_36 <= nl_res_rsci_d_53_36[17:0];
      res_rsci_d_521_504 <= nl_res_rsci_d_521_504[17:0];
      res_rsci_d_71_54 <= nl_res_rsci_d_71_54[17:0];
      res_rsci_d_503_486 <= nl_res_rsci_d_503_486[17:0];
      res_rsci_d_89_72 <= nl_res_rsci_d_89_72[17:0];
      res_rsci_d_485_468 <= nl_res_rsci_d_485_468[17:0];
      res_rsci_d_107_90 <= nl_res_rsci_d_107_90[17:0];
      res_rsci_d_467_450 <= nl_res_rsci_d_467_450[17:0];
      res_rsci_d_125_108 <= nl_res_rsci_d_125_108[17:0];
      res_rsci_d_449_432 <= nl_res_rsci_d_449_432[17:0];
      res_rsci_d_143_126 <= nl_res_rsci_d_143_126[17:0];
      res_rsci_d_431_414 <= nl_res_rsci_d_431_414[17:0];
      res_rsci_d_161_144 <= nl_res_rsci_d_161_144[17:0];
      res_rsci_d_413_396 <= nl_res_rsci_d_413_396[17:0];
      res_rsci_d_179_162 <= nl_res_rsci_d_179_162[17:0];
      res_rsci_d_395_378 <= nl_res_rsci_d_395_378[17:0];
      res_rsci_d_197_180 <= nl_res_rsci_d_197_180[17:0];
      res_rsci_d_377_360 <= nl_res_rsci_d_377_360[17:0];
      res_rsci_d_215_198 <= nl_res_rsci_d_215_198[17:0];
      res_rsci_d_359_342 <= nl_res_rsci_d_359_342[17:0];
      res_rsci_d_233_216 <= nl_res_rsci_d_233_216[17:0];
      res_rsci_d_341_324 <= nl_res_rsci_d_341_324[17:0];
      res_rsci_d_251_234 <= nl_res_rsci_d_251_234[17:0];
      res_rsci_d_323_306 <= nl_res_rsci_d_323_306[17:0];
      res_rsci_d_269_252 <= nl_res_rsci_d_269_252[17:0];
      res_rsci_d_305_288 <= nl_res_rsci_d_305_288[17:0];
      res_rsci_d_287_270 <= nl_res_rsci_d_287_270[17:0];
    end
  end
  assign nl_Result_acc_94_nl = conv_s2s_25_26({(~ (data_rsci_idat[161:144])) , 7'b0000001})
      + conv_s2s_19_26({Result_Result_conc_52_18_10 , (~ (data_rsci_idat[153:144]))});
  assign Result_acc_94_nl = nl_Result_acc_94_nl[25:0];
  assign nl_Result_acc_242_nl = conv_s2u_19_21(readslicef_26_19_7((Result_acc_94_nl)))
      + ({(~ (data_rsci_idat[161:144])) , 3'b001});
  assign Result_acc_242_nl = nl_Result_acc_242_nl[20:0];
  assign nl_Result_acc_87_nl = ({(~ (data_rsci_idat[35:18])) , 5'b00000}) + conv_s2s_21_23(MultLoop_acc_759_sdt_1);
  assign Result_acc_87_nl = nl_Result_acc_87_nl[22:0];
  assign nl_Result_acc_70_nl = conv_s2s_23_25(Result_acc_87_nl) + ({(data_rsci_idat[35:18])
      , 7'b0100000});
  assign Result_acc_70_nl = nl_Result_acc_70_nl[24:0];
  assign nl_Result_acc_90_nl = ({(data_rsci_idat[89:72]) , 6'b010000}) + conv_s2s_22_24({(~
      (data_rsci_idat[89:72])) , 4'b0001}) + conv_s2s_19_24({Result_Result_conc_54_18_8
      , (~ (data_rsci_idat[79:72]))});
  assign Result_acc_90_nl = nl_Result_acc_90_nl[23:0];
  assign nl_Result_acc_244_nl = conv_s2u_16_18(readslicef_24_16_8((Result_acc_90_nl)))
      + (~ (data_rsci_idat[89:72]));
  assign Result_acc_244_nl = nl_Result_acc_244_nl[17:0];
  assign nl_MultLoop_acc_416_nl = conv_s2s_16_17(readslicef_25_16_9((Result_acc_70_nl)))
      + conv_s2s_16_17(readslicef_18_16_2((Result_acc_244_nl)));
  assign MultLoop_acc_416_nl = nl_MultLoop_acc_416_nl[16:0];
  assign nl_MultLoop_acc_419_nl = (readslicef_21_18_3((Result_acc_242_nl))) + conv_s2s_17_18(MultLoop_acc_416_nl);
  assign MultLoop_acc_419_nl = nl_MultLoop_acc_419_nl[17:0];
  assign nl_MultLoop_acc_1347_nl = conv_s2s_8_9(Result_acc_71_itm_17_7[10:3]) + 9'b111111101;
  assign MultLoop_acc_1347_nl = nl_MultLoop_acc_1347_nl[8:0];
  assign nl_MultLoop_acc_414_nl = MultLoop_acc_1350_itm_18_5 + conv_s2s_12_14({(MultLoop_acc_1347_nl)
      , (Result_acc_71_itm_17_7[2:0])});
  assign MultLoop_acc_414_nl = nl_MultLoop_acc_414_nl[13:0];
  assign nl_MultLoop_acc_415_nl = MultLoop_acc_1348_itm_18_3 + conv_s2s_14_16(MultLoop_acc_414_nl);
  assign MultLoop_acc_415_nl = nl_MultLoop_acc_415_nl[15:0];
  assign nl_MultLoop_acc_418_nl = conv_s2s_16_17(MultLoop_acc_415_nl) + MultLoop_acc_353_itm_22_6;
  assign MultLoop_acc_418_nl = nl_MultLoop_acc_418_nl[16:0];
  assign nl_MultLoop_acc_421_nl = (MultLoop_acc_419_nl) + conv_s2s_17_18(MultLoop_acc_418_nl);
  assign MultLoop_acc_421_nl = nl_MultLoop_acc_421_nl[17:0];
  assign nl_Result_acc_92_nl = ({(data_rsci_idat[143:126]) , 4'b0001}) + conv_s2s_19_22({Result_Result_conc_48_18_9
      , (~ (data_rsci_idat[134:126]))});
  assign Result_acc_92_nl = nl_Result_acc_92_nl[21:0];
  assign nl_Result_acc_246_nl = conv_s2u_13_18(readslicef_22_13_9((Result_acc_92_nl)))
      + (~ (data_rsci_idat[143:126]));
  assign Result_acc_246_nl = nl_Result_acc_246_nl[17:0];
  assign nl_Result_acc_85_nl = (~ (data_rsci_idat[17:0])) + conv_s2s_15_18({MultLoop_acc_1254_cse_1
      , (data_rsci_idat[6:4])});
  assign Result_acc_85_nl = nl_Result_acc_85_nl[17:0];
  assign nl_Result_acc_79_nl = conv_s2u_18_22(Result_acc_85_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[17:0])) , 3'b001});
  assign Result_acc_79_nl = nl_Result_acc_79_nl[21:0];
  assign nl_MultLoop_acc_417_nl = conv_s2s_17_18(readslicef_18_17_1((Result_acc_246_nl)))
      + conv_s2s_16_18(readslicef_22_16_6((Result_acc_79_nl)));
  assign MultLoop_acc_417_nl = nl_MultLoop_acc_417_nl[17:0];
  assign nl_MultLoop_acc_420_nl = (MultLoop_acc_417_nl) + (~ (data_rsci_idat[125:108]));
  assign MultLoop_acc_420_nl = nl_MultLoop_acc_420_nl[17:0];
  assign nl_res_rsci_d_575_558  = (MultLoop_acc_421_nl) + (MultLoop_acc_420_nl);
  assign nl_MultLoop_acc_1136_nl = conv_s2s_18_19(data_rsci_idat[71:54]) + conv_s2s_14_19({MultLoop_acc_1213_cse_1
      , (data_rsci_idat[63:59])});
  assign MultLoop_acc_1136_nl = nl_MultLoop_acc_1136_nl[18:0];
  assign nl_MultLoop_acc_16_nl = conv_s2u_19_23(MultLoop_acc_1136_nl) + ({(~ (data_rsci_idat[71:54]))
      , 5'b00000});
  assign MultLoop_acc_16_nl = nl_MultLoop_acc_16_nl[22:0];
  assign nl_MultLoop_acc_294_nl = conv_s2u_15_19(data_rsci_idat[143:129]) + conv_s2u_18_19(data_rsci_idat[143:126]);
  assign MultLoop_acc_294_nl = nl_MultLoop_acc_294_nl[18:0];
  assign nl_MultLoop_acc_1144_nl = (readslicef_23_18_5((MultLoop_acc_16_nl))) + (readslicef_19_18_1((MultLoop_acc_294_nl)));
  assign MultLoop_acc_1144_nl = nl_MultLoop_acc_1144_nl[17:0];
  assign nl_MultLoop_acc_12_nl = conv_s2s_18_22(~ (data_rsci_idat[17:0])) + ({(data_rsci_idat[17:0])
      , 4'b0001});
  assign MultLoop_acc_12_nl = nl_MultLoop_acc_12_nl[21:0];
  assign nl_MultLoop_acc_18_nl = conv_s2s_18_20(~ (data_rsci_idat[107:90])) + ({(data_rsci_idat[107:90])
      , 2'b01});
  assign MultLoop_acc_18_nl = nl_MultLoop_acc_18_nl[19:0];
  assign nl_MultLoop_acc_1343_nl = conv_s2u_9_10(data_rsci_idat[161:153]) + 10'b0110101111;
  assign MultLoop_acc_1343_nl = nl_MultLoop_acc_1343_nl[9:0];
  assign nl_MultLoop_acc_1138_nl = conv_s2s_13_14(readslicef_20_13_7((MultLoop_acc_18_nl)))
      + conv_u2s_11_14({(MultLoop_acc_1343_nl) , (data_rsci_idat[152])});
  assign MultLoop_acc_1138_nl = nl_MultLoop_acc_1138_nl[13:0];
  assign nl_MultLoop_acc_1124_nl = (~ (data_rsci_idat[89:72])) + conv_s2s_15_18(data_rsci_idat[89:75]);
  assign MultLoop_acc_1124_nl = nl_MultLoop_acc_1124_nl[17:0];
  assign nl_MultLoop_acc_293_nl = conv_s2u_18_20(MultLoop_acc_1124_nl) + ({(data_rsci_idat[89:72])
      , 2'b01});
  assign MultLoop_acc_293_nl = nl_MultLoop_acc_293_nl[19:0];
  assign nl_MultLoop_acc_1143_nl = (data_rsci_idat[161:144]) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_12_nl)))
      + conv_s2s_14_18(MultLoop_acc_1138_nl) + conv_s2s_14_18(MultLoop_acc_19_itm_19_3[16:3])
      + conv_s2s_14_18(readslicef_20_14_6((MultLoop_acc_293_nl)));
  assign MultLoop_acc_1143_nl = nl_MultLoop_acc_1143_nl[17:0];
  assign nl_MultLoop_acc_1146_nl = (MultLoop_acc_1144_nl) + (MultLoop_acc_1143_nl);
  assign MultLoop_acc_1146_nl = nl_MultLoop_acc_1146_nl[17:0];
  assign nl_MultLoop_acc_1127_nl = conv_s2s_20_21({(data_rsci_idat[179:162]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[179:162]) + conv_s2s_15_21({MultLoop_acc_1273_cse_1
      , (data_rsci_idat[170:166])});
  assign MultLoop_acc_1127_nl = nl_MultLoop_acc_1127_nl[20:0];
  assign nl_MultLoop_acc_22_nl = conv_s2u_21_23(MultLoop_acc_1127_nl) + ({(~ (data_rsci_idat[179:162]))
      , 5'b00000});
  assign MultLoop_acc_22_nl = nl_MultLoop_acc_22_nl[22:0];
  assign nl_MultLoop_acc_1129_nl = ({(~ (data_rsci_idat[35:18])) , 2'b00}) + conv_s2s_19_20(MultLoop_acc_875_cse_1);
  assign MultLoop_acc_1129_nl = nl_MultLoop_acc_1129_nl[19:0];
  assign nl_MultLoop_acc_292_nl = conv_s2u_20_25(MultLoop_acc_1129_nl) + ({(data_rsci_idat[35:18])
      , 7'b0000100});
  assign MultLoop_acc_292_nl = nl_MultLoop_acc_292_nl[24:0];
  assign nl_MultLoop_acc_1142_nl = conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_22_nl)))
      + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_292_nl)));
  assign MultLoop_acc_1142_nl = nl_MultLoop_acc_1142_nl[17:0];
  assign nl_MultLoop_acc_1131_nl = ({(data_rsci_idat[53:36]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_214_18_10
      , (~ (data_rsci_idat[45:36]))});
  assign MultLoop_acc_1131_nl = nl_MultLoop_acc_1131_nl[19:0];
  assign nl_MultLoop_acc_1132_nl = ({(~ (data_rsci_idat[53:36])) , 4'b0000}) + conv_s2s_20_22(MultLoop_acc_1131_nl);
  assign MultLoop_acc_1132_nl = nl_MultLoop_acc_1132_nl[21:0];
  assign nl_MultLoop_acc_1134_nl = conv_s2s_26_27({(~ (data_rsci_idat[53:36])) ,
      8'b01000000}) + conv_s2s_24_27({(~ (data_rsci_idat[53:36])) , 6'b010000}) +
      conv_s2s_22_27(MultLoop_acc_1132_nl);
  assign MultLoop_acc_1134_nl = nl_MultLoop_acc_1134_nl[26:0];
  assign nl_MultLoop_acc_1346_nl = conv_s2u_19_20(readslicef_27_19_8((MultLoop_acc_1134_nl)))
      + ({(~ (data_rsci_idat[53:36])) , 2'b01});
  assign MultLoop_acc_1346_nl = nl_MultLoop_acc_1346_nl[19:0];
  assign nl_MultLoop_acc_1145_nl = (MultLoop_acc_1142_nl) + (readslicef_20_18_2((MultLoop_acc_1346_nl)));
  assign MultLoop_acc_1145_nl = nl_MultLoop_acc_1145_nl[17:0];
  assign nl_res_rsci_d_17_0  = (MultLoop_acc_1146_nl) + (MultLoop_acc_1145_nl);
  assign nl_Result_acc_236_nl = conv_s2s_9_10(data_rsci_idat[35:27]) + 10'b0000000001;
  assign Result_acc_236_nl = nl_Result_acc_236_nl[9:0];
  assign nl_Result_acc_106_nl = (~ (data_rsci_idat[35:18])) + conv_s2s_17_18({(Result_acc_236_nl)
      , (data_rsci_idat[26:20])});
  assign Result_acc_106_nl = nl_Result_acc_106_nl[17:0];
  assign nl_Result_acc_107_nl = ({(data_rsci_idat[35:18]) , 2'b01}) + conv_s2s_18_20(Result_acc_106_nl);
  assign Result_acc_107_nl = nl_Result_acc_107_nl[19:0];
  assign nl_Result_acc_108_nl = conv_s2s_22_23({(data_rsci_idat[35:18]) , 4'b0000})
      + conv_s2s_20_23(Result_acc_107_nl);
  assign Result_acc_108_nl = nl_Result_acc_108_nl[22:0];
  assign nl_Result_acc_237_nl = conv_s2u_16_18(readslicef_23_16_7((Result_acc_108_nl)))
      + (~ (data_rsci_idat[35:18]));
  assign Result_acc_237_nl = nl_Result_acc_237_nl[17:0];
  assign nl_Result_acc_60_nl = conv_s2s_18_27(~ (data_rsci_idat[89:72])) + ({(data_rsci_idat[89:72])
      , 9'b000000001});
  assign Result_acc_60_nl = nl_Result_acc_60_nl[26:0];
  assign nl_Result_acc_110_nl = ({(data_rsci_idat[107:90]) , 2'b01}) + conv_s2s_19_20({Result_Result_conc_58_18_9
      , (~ (data_rsci_idat[98:90]))});
  assign Result_acc_110_nl = nl_Result_acc_110_nl[19:0];
  assign nl_Result_acc_239_nl = conv_s2u_11_18(readslicef_20_11_9((Result_acc_110_nl)))
      + (~ (data_rsci_idat[107:90]));
  assign Result_acc_239_nl = nl_Result_acc_239_nl[17:0];
  assign nl_Result_acc_240_nl =  -conv_s2s_11_12(data_rsci_idat[143:133]);
  assign Result_acc_240_nl = nl_Result_acc_240_nl[11:0];
  assign nl_Result_acc_63_nl = conv_s2s_25_26({(~ (data_rsci_idat[143:126])) , 7'b0010000})
      + conv_s2s_22_26({(~ (data_rsci_idat[143:126])) , 4'b0100}) + conv_s2s_20_26({(~
      (data_rsci_idat[143:126])) , 2'b01}) + conv_s2s_19_26({(Result_acc_240_nl)
      , (~ (data_rsci_idat[132:126]))});
  assign Result_acc_63_nl = nl_Result_acc_63_nl[25:0];
  assign nl_MultLoop_acc_429_nl = conv_s2s_17_18(readslicef_18_17_1((Result_acc_237_nl)))
      + conv_s2s_17_18(readslicef_27_17_10((Result_acc_60_nl))) + conv_s2s_17_18(readslicef_18_17_1((Result_acc_239_nl)))
      + conv_s2s_17_18(readslicef_26_17_9((Result_acc_63_nl)));
  assign MultLoop_acc_429_nl = nl_MultLoop_acc_429_nl[17:0];
  assign nl_Result_acc_115_nl = conv_s2s_23_24({(~ (data_rsci_idat[161:144])) , 5'b01000})
      + conv_s2s_21_24({(~ (data_rsci_idat[161:144])) , 3'b001}) + conv_s2s_18_24(~
      (data_rsci_idat[161:144]));
  assign Result_acc_115_nl = nl_Result_acc_115_nl[23:0];
  assign nl_Result_acc_64_nl = conv_s2s_24_27(Result_acc_115_nl) + ({(data_rsci_idat[161:144])
      , 9'b000100000});
  assign Result_acc_64_nl = nl_Result_acc_64_nl[26:0];
  assign nl_Result_acc_96_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_14_18({Result_Result_conc_50_13_2
      , (data_rsci_idat[42:41])});
  assign Result_acc_96_nl = nl_Result_acc_96_nl[17:0];
  assign nl_Result_acc_66_nl = conv_s2u_18_21(Result_acc_96_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[53:36])) , 2'b01});
  assign Result_acc_66_nl = nl_Result_acc_66_nl[20:0];
  assign nl_MultLoop_acc_424_nl = conv_s2s_17_18(readslicef_27_17_10((Result_acc_64_nl)))
      + conv_s2s_16_18(readslicef_21_16_5((Result_acc_66_nl)));
  assign MultLoop_acc_424_nl = nl_MultLoop_acc_424_nl[17:0];
  assign nl_Result_acc_248_nl = ({(data_rsci_idat[17:0]) , 2'b01}) + conv_s2u_19_20(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_5_cse_1[21:3]);
  assign Result_acc_248_nl = nl_Result_acc_248_nl[19:0];
  assign nl_Result_acc_232_nl = conv_s2u_16_19(readslicef_20_16_4((Result_acc_248_nl)))
      + conv_s2u_18_19(data_rsci_idat[17:0]);
  assign Result_acc_232_nl = nl_Result_acc_232_nl[18:0];
  assign nl_MultLoop_acc_428_nl = (MultLoop_acc_424_nl) + (readslicef_19_18_1((Result_acc_232_nl)));
  assign MultLoop_acc_428_nl = nl_MultLoop_acc_428_nl[17:0];
  assign nl_Result_acc_104_nl = conv_s2s_20_21({(~ (data_rsci_idat[179:162])) , 2'b01})
      + conv_s2s_18_21(MultLoop_acc_634_cse_1);
  assign Result_acc_104_nl = nl_Result_acc_104_nl[20:0];
  assign nl_Result_acc_68_nl = conv_s2u_21_23(Result_acc_104_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[179:162])) , 4'b0100});
  assign Result_acc_68_nl = nl_Result_acc_68_nl[22:0];
  assign nl_MultLoop_acc_422_nl = conv_s2s_16_17(readslicef_23_16_7((Result_acc_68_nl)))
      + 17'b00000001000000111;
  assign MultLoop_acc_422_nl = nl_MultLoop_acc_422_nl[16:0];
  assign nl_Result_acc_98_nl = (~ (data_rsci_idat[71:54])) + conv_s2s_14_18({MultLoop_acc_1148_cse_1
      , (data_rsci_idat[60:59])});
  assign Result_acc_98_nl = nl_Result_acc_98_nl[17:0];
  assign nl_Result_acc_67_nl = conv_s2u_18_21(Result_acc_98_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[71:54])) , 2'b01});
  assign Result_acc_67_nl = nl_Result_acc_67_nl[20:0];
  assign nl_Result_acc_234_nl = conv_s2s_12_13(data_rsci_idat[125:114]) + 13'b0000000000001;
  assign Result_acc_234_nl = nl_Result_acc_234_nl[12:0];
  assign nl_Result_acc_101_nl = conv_s2s_20_21({(data_rsci_idat[125:108]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[125:108]) + conv_s2s_17_21({(Result_acc_234_nl)
      , (data_rsci_idat[113:110])});
  assign Result_acc_101_nl = nl_Result_acc_101_nl[20:0];
  assign nl_Result_acc_62_nl = conv_s2u_21_22(Result_acc_101_nl) + ({(~ (data_rsci_idat[125:108]))
      , 4'b0000});
  assign Result_acc_62_nl = nl_Result_acc_62_nl[21:0];
  assign nl_res_rsci_d_557_540  = (MultLoop_acc_429_nl) + (MultLoop_acc_428_nl) +
      conv_s2s_17_18(MultLoop_acc_422_nl) + conv_s2s_16_18(readslicef_21_16_5((Result_acc_67_nl)))
      + conv_s2s_16_18(readslicef_22_16_6((Result_acc_62_nl)));
  assign nl_MultLoop_acc_1330_nl = conv_s2u_16_19(MultLoop_acc_213_itm_22_7) + conv_s2u_18_19(data_rsci_idat[143:126]);
  assign MultLoop_acc_1330_nl = nl_MultLoop_acc_1330_nl[18:0];
  assign nl_MultLoop_acc_1098_nl = conv_s2s_18_19(data_rsci_idat[89:72]) + conv_s2s_13_19(data_rsci_idat[89:77]);
  assign MultLoop_acc_1098_nl = nl_MultLoop_acc_1098_nl[18:0];
  assign nl_MultLoop_acc_296_nl = conv_s2u_19_21(MultLoop_acc_1098_nl) + conv_s2u_20_21({(data_rsci_idat[89:72])
      , 2'b00});
  assign MultLoop_acc_296_nl = nl_MultLoop_acc_296_nl[20:0];
  assign nl_MultLoop_acc_1331_nl =  -conv_s2s_10_11(data_rsci_idat[107:98]);
  assign MultLoop_acc_1331_nl = nl_MultLoop_acc_1331_nl[10:0];
  assign nl_MultLoop_acc_1100_nl = ({(data_rsci_idat[107:90]) , 4'b0001}) + conv_s2s_19_22({(MultLoop_acc_1331_nl)
      , (~ (data_rsci_idat[97:90]))});
  assign MultLoop_acc_1100_nl = nl_MultLoop_acc_1100_nl[21:0];
  assign nl_MultLoop_acc_1101_nl = conv_s2s_24_25({(data_rsci_idat[107:90]) , 6'b000000})
      + conv_s2s_22_25(MultLoop_acc_1100_nl);
  assign MultLoop_acc_1101_nl = nl_MultLoop_acc_1101_nl[24:0];
  assign nl_MultLoop_acc_1332_nl = conv_s2u_17_18(readslicef_25_17_8((MultLoop_acc_1101_nl)))
      + (~ (data_rsci_idat[107:90]));
  assign MultLoop_acc_1332_nl = nl_MultLoop_acc_1332_nl[17:0];
  assign nl_MultLoop_acc_1333_nl =  -conv_s2s_10_11(data_rsci_idat[17:8]);
  assign MultLoop_acc_1333_nl = nl_MultLoop_acc_1333_nl[10:0];
  assign nl_MultLoop_acc_1093_nl = ({(data_rsci_idat[17:0]) , 6'b000001}) + conv_s2s_19_24({(MultLoop_acc_1333_nl)
      , (~ (data_rsci_idat[7:0]))});
  assign MultLoop_acc_1093_nl = nl_MultLoop_acc_1093_nl[23:0];
  assign nl_MultLoop_acc_1334_nl = conv_s2u_16_18(readslicef_24_16_8((MultLoop_acc_1093_nl)))
      + (~ (data_rsci_idat[17:0]));
  assign MultLoop_acc_1334_nl = nl_MultLoop_acc_1334_nl[17:0];
  assign nl_MultLoop_acc_1115_nl = (readslicef_18_16_2((MultLoop_acc_1334_nl))) +
      16'b0000001100101001;
  assign MultLoop_acc_1115_nl = nl_MultLoop_acc_1115_nl[15:0];
  assign nl_MultLoop_acc_1121_nl = conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_1330_nl)))
      + conv_s2s_17_18(readslicef_21_17_4((MultLoop_acc_296_nl))) + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_1332_nl)))
      + conv_s2s_16_18(MultLoop_acc_1115_nl);
  assign MultLoop_acc_1121_nl = nl_MultLoop_acc_1121_nl[17:0];
  assign nl_MultLoop_acc_1103_nl = conv_s2s_24_25({(~ (data_rsci_idat[35:18])) ,
      6'b001000}) + conv_s2s_22_25(MultLoop_acc_839_cse_1);
  assign MultLoop_acc_1103_nl = nl_MultLoop_acc_1103_nl[24:0];
  assign nl_MultLoop_acc_24_nl = conv_s2s_25_28(MultLoop_acc_1103_nl) + ({(data_rsci_idat[35:18])
      , 10'b0001000000});
  assign MultLoop_acc_24_nl = nl_MultLoop_acc_24_nl[27:0];
  assign nl_MultLoop_acc_1106_nl = ({(data_rsci_idat[53:36]) , 5'b00100}) + conv_s2s_20_23({(~
      (data_rsci_idat[53:36])) , 2'b01}) + conv_s2s_19_23({MultLoop_MultLoop_conc_214_18_10
      , (~ (data_rsci_idat[45:36]))});
  assign MultLoop_acc_1106_nl = nl_MultLoop_acc_1106_nl[22:0];
  assign nl_MultLoop_acc_1336_nl = conv_s2u_18_19(data_rsci_idat[53:36]) + conv_s2u_15_19(readslicef_23_15_8((MultLoop_acc_1106_nl)));
  assign MultLoop_acc_1336_nl = nl_MultLoop_acc_1336_nl[18:0];
  assign nl_MultLoop_acc_1337_nl = conv_s2u_17_18(readslicef_19_17_2((MultLoop_acc_1336_nl)))
      + (~ (data_rsci_idat[53:36]));
  assign MultLoop_acc_1337_nl = nl_MultLoop_acc_1337_nl[17:0];
  assign nl_MultLoop_acc_1120_nl = (readslicef_28_18_10((MultLoop_acc_24_nl))) +
      (MultLoop_acc_1337_nl);
  assign MultLoop_acc_1120_nl = nl_MultLoop_acc_1120_nl[17:0];
  assign nl_MultLoop_acc_1123_nl = (MultLoop_acc_1121_nl) + (MultLoop_acc_1120_nl);
  assign MultLoop_acc_1123_nl = nl_MultLoop_acc_1123_nl[17:0];
  assign nl_MultLoop_acc_1338_nl = conv_s2s_10_11(data_rsci_idat[71:62]) + 11'b00000000001;
  assign MultLoop_acc_1338_nl = nl_MultLoop_acc_1338_nl[10:0];
  assign nl_MultLoop_acc_1110_nl = conv_s2s_22_23({(data_rsci_idat[71:54]) , 4'b0000})
      + conv_s2s_18_23(data_rsci_idat[71:54]) + conv_s2s_17_23({(MultLoop_acc_1338_nl)
      , (data_rsci_idat[61:56])});
  assign MultLoop_acc_1110_nl = nl_MultLoop_acc_1110_nl[22:0];
  assign nl_MultLoop_acc_1339_nl = conv_s2u_17_18(readslicef_23_17_6((MultLoop_acc_1110_nl)))
      + (~ (data_rsci_idat[71:54]));
  assign MultLoop_acc_1339_nl = nl_MultLoop_acc_1339_nl[17:0];
  assign nl_MultLoop_acc_1111_nl = ({(data_rsci_idat[125:108]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[125:108]));
  assign MultLoop_acc_1111_nl = nl_MultLoop_acc_1111_nl[20:0];
  assign nl_MultLoop_acc_29_nl = conv_s2s_21_24(MultLoop_acc_1111_nl) + conv_s2s_23_24({(data_rsci_idat[125:108])
      , 5'b00000});
  assign MultLoop_acc_29_nl = nl_MultLoop_acc_29_nl[23:0];
  assign nl_MultLoop_acc_1119_nl = (MultLoop_acc_1339_nl) + (readslicef_24_18_6((MultLoop_acc_29_nl)));
  assign MultLoop_acc_1119_nl = nl_MultLoop_acc_1119_nl[17:0];
  assign nl_MultLoop_acc_1113_nl = (~ (data_rsci_idat[179:162])) + conv_s2s_17_18({MultLoop_acc_1273_cse_1
      , (data_rsci_idat[170:164])});
  assign MultLoop_acc_1113_nl = nl_MultLoop_acc_1113_nl[17:0];
  assign nl_MultLoop_acc_1114_nl = conv_s2s_20_21({(~ (data_rsci_idat[179:162]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_1113_nl);
  assign MultLoop_acc_1114_nl = nl_MultLoop_acc_1114_nl[20:0];
  assign nl_MultLoop_acc_297_nl = conv_s2u_21_26(MultLoop_acc_1114_nl) + conv_s2u_25_26({(~
      (data_rsci_idat[179:162])) , 7'b0000100});
  assign MultLoop_acc_297_nl = nl_MultLoop_acc_297_nl[25:0];
  assign nl_MultLoop_acc_1095_nl = ({(~ (data_rsci_idat[161:144])) , 5'b00000}) +
      conv_s2s_20_23(MultLoop_acc_892_cse_1);
  assign MultLoop_acc_1095_nl = nl_MultLoop_acc_1095_nl[22:0];
  assign nl_MultLoop_acc_1096_nl = conv_s2s_25_26({(~ (data_rsci_idat[161:144]))
      , 7'b0100000}) + conv_s2s_23_26(MultLoop_acc_1095_nl);
  assign MultLoop_acc_1096_nl = nl_MultLoop_acc_1096_nl[25:0];
  assign nl_MultLoop_acc_1341_nl = conv_s2u_19_20(readslicef_26_19_7((MultLoop_acc_1096_nl)))
      + ({(data_rsci_idat[161:144]) , 2'b01});
  assign MultLoop_acc_1341_nl = nl_MultLoop_acc_1341_nl[19:0];
  assign nl_MultLoop_acc_1118_nl = (readslicef_26_18_8((MultLoop_acc_297_nl))) +
      conv_s2s_17_18(readslicef_20_17_3((MultLoop_acc_1341_nl)));
  assign MultLoop_acc_1118_nl = nl_MultLoop_acc_1118_nl[17:0];
  assign nl_MultLoop_acc_1122_nl = (MultLoop_acc_1119_nl) + (MultLoop_acc_1118_nl);
  assign MultLoop_acc_1122_nl = nl_MultLoop_acc_1122_nl[17:0];
  assign nl_res_rsci_d_35_18  = (MultLoop_acc_1123_nl) + (MultLoop_acc_1122_nl);
  assign nl_Result_acc_223_nl = conv_s2s_12_13(data_rsci_idat[143:132]) + 13'b0000000000001;
  assign Result_acc_223_nl = nl_Result_acc_223_nl[12:0];
  assign nl_Result_acc_128_nl = (~ (data_rsci_idat[143:126])) + conv_s2s_16_18({(Result_acc_223_nl)
      , (data_rsci_idat[131:129])});
  assign Result_acc_128_nl = nl_Result_acc_128_nl[17:0];
  assign nl_Result_acc_55_nl = conv_s2u_18_22(Result_acc_128_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[143:126])) , 3'b001});
  assign Result_acc_55_nl = nl_Result_acc_55_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_15_nl = conv_s2u_16_19(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_4_itm_18_2_1[16:1])
      + conv_s2u_18_19(data_rsci_idat[17:0]);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_15_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_15_nl[18:0];
  assign nl_MultLoop_acc_433_nl = (readslicef_22_17_5((Result_acc_55_nl))) + conv_s2s_16_17(readslicef_19_16_3((nnet_product_input_t_config2_weight_t_config2_accum_t_acc_15_nl)));
  assign MultLoop_acc_433_nl = nl_MultLoop_acc_433_nl[16:0];
  assign nl_Result_acc_224_nl =  -conv_s2s_9_10(data_rsci_idat[35:27]);
  assign Result_acc_224_nl = nl_Result_acc_224_nl[9:0];
  assign nl_Result_acc_130_nl = ({(data_rsci_idat[35:18]) , 5'b00001}) + conv_s2s_19_23({(Result_acc_224_nl)
      , (~ (data_rsci_idat[26:18]))});
  assign Result_acc_130_nl = nl_Result_acc_130_nl[22:0];
  assign nl_Result_acc_225_nl = (~ (data_rsci_idat[35:18])) + conv_s2s_16_18(readslicef_23_16_7((Result_acc_130_nl)));
  assign Result_acc_225_nl = nl_Result_acc_225_nl[17:0];
  assign nl_Result_acc_226_nl = conv_s2u_18_21(Result_acc_225_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[35:18])) , 2'b01});
  assign Result_acc_226_nl = nl_Result_acc_226_nl[20:0];
  assign nl_MultLoop_acc_437_nl = conv_s2s_17_18(MultLoop_acc_433_nl) + (readslicef_21_18_3((Result_acc_226_nl)));
  assign MultLoop_acc_437_nl = nl_MultLoop_acc_437_nl[17:0];
  assign nl_Result_acc_47_nl = conv_s2s_26_27({(~ (data_rsci_idat[71:54])) , 8'b00100000})
      + conv_s2s_23_27({(~ (data_rsci_idat[71:54])) , 5'b00100}) + conv_s2s_20_27({(~
      (data_rsci_idat[71:54])) , 2'b01}) + conv_s2s_19_27({Result_Result_conc_64_18_8
      , (~ (data_rsci_idat[61:54]))});
  assign Result_acc_47_nl = nl_Result_acc_47_nl[26:0];
  assign nl_Result_acc_251_nl = conv_s2u_19_22(MultLoop_acc_1390_itm_22_4_1) + ({(data_rsci_idat[161:144])
      , 4'b0001});
  assign Result_acc_251_nl = nl_Result_acc_251_nl[21:0];
  assign nl_MultLoop_acc_436_nl = (readslicef_27_18_9((Result_acc_47_nl))) + (readslicef_22_18_4((Result_acc_251_nl)));
  assign MultLoop_acc_436_nl = nl_MultLoop_acc_436_nl[17:0];
  assign nl_MultLoop_acc_439_nl = (MultLoop_acc_437_nl) + (MultLoop_acc_436_nl);
  assign MultLoop_acc_439_nl = nl_MultLoop_acc_439_nl[17:0];
  assign nl_Result_acc_120_nl = ({(~ (data_rsci_idat[89:72])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[89:72])
      + conv_s2s_15_20(data_rsci_idat[89:75]);
  assign Result_acc_120_nl = nl_Result_acc_120_nl[19:0];
  assign nl_Result_acc_121_nl = conv_s2s_22_23({(~ (data_rsci_idat[89:72])) , 4'b0100})
      + conv_s2s_20_23(Result_acc_120_nl);
  assign Result_acc_121_nl = nl_Result_acc_121_nl[22:0];
  assign nl_Result_acc_54_nl = conv_s2u_23_24(Result_acc_121_nl) + ({(data_rsci_idat[89:72])
      , 6'b010000});
  assign Result_acc_54_nl = nl_Result_acc_54_nl[23:0];
  assign nl_Result_acc_118_nl = conv_s2s_20_21({(~ (data_rsci_idat[179:162])) , 2'b01})
      + conv_s2s_18_21(~ (data_rsci_idat[179:162]));
  assign Result_acc_118_nl = nl_Result_acc_118_nl[20:0];
  assign nl_Result_acc_53_nl = conv_s2s_21_23(Result_acc_118_nl) + ({(data_rsci_idat[179:162])
      , 5'b00100});
  assign Result_acc_53_nl = nl_Result_acc_53_nl[22:0];
  assign nl_MultLoop_acc_1329_nl = conv_s2s_12_13(Result_acc_46_itm_17_4[13:2]) +
      13'b0000001000101;
  assign MultLoop_acc_1329_nl = nl_MultLoop_acc_1329_nl[12:0];
  assign nl_Result_acc_49_nl = conv_s2s_25_26({(~ (data_rsci_idat[107:90])) , 7'b0100000})
      + conv_s2s_23_26({(~ (data_rsci_idat[107:90])) , 5'b00100}) + conv_s2s_20_26({(~
      (data_rsci_idat[107:90])) , 2'b01}) + conv_s2s_19_26({Result_Result_conc_60_18_7
      , (~ (data_rsci_idat[96:90]))});
  assign Result_acc_49_nl = nl_Result_acc_49_nl[25:0];
  assign nl_Result_acc_229_nl =  -conv_s2s_10_11(data_rsci_idat[125:116]);
  assign Result_acc_229_nl = nl_Result_acc_229_nl[10:0];
  assign nl_Result_acc_126_nl = ({(data_rsci_idat[125:108]) , 4'b0001}) + conv_s2s_19_22({(Result_acc_229_nl)
      , (~ (data_rsci_idat[115:108]))});
  assign Result_acc_126_nl = nl_Result_acc_126_nl[21:0];
  assign nl_Result_acc_230_nl = conv_s2u_14_18(readslicef_22_14_8((Result_acc_126_nl)))
      + (~ (data_rsci_idat[125:108]));
  assign Result_acc_230_nl = nl_Result_acc_230_nl[17:0];
  assign nl_res_rsci_d_539_522  = (MultLoop_acc_439_nl) + conv_s2s_17_18(readslicef_24_17_7((Result_acc_54_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((Result_acc_53_nl))) + conv_s2s_15_18({(MultLoop_acc_1329_nl)
      , (Result_acc_46_itm_17_4[1:0])}) + conv_s2s_17_18(readslicef_26_17_9((Result_acc_49_nl)))
      + conv_s2s_17_18(readslicef_18_17_1((Result_acc_230_nl)));
  assign nl_MultLoop_acc_1078_nl = ({(data_rsci_idat[107:90]) , 7'b0100000}) + conv_s2s_23_25({(~
      (data_rsci_idat[107:90])) , 5'b01000}) + conv_s2s_21_25({(~ (data_rsci_idat[107:90]))
      , 3'b001}) + conv_s2s_19_25({Result_Result_conc_58_18_9 , (~ (data_rsci_idat[98:90]))});
  assign MultLoop_acc_1078_nl = nl_MultLoop_acc_1078_nl[24:0];
  assign nl_MultLoop_acc_1324_nl = conv_s2u_16_18(readslicef_25_16_9((MultLoop_acc_1078_nl)))
      + (~ (data_rsci_idat[107:90]));
  assign MultLoop_acc_1324_nl = nl_MultLoop_acc_1324_nl[17:0];
  assign nl_MultLoop_acc_1385_nl = conv_s2u_16_19(MultLoop_acc_123_itm_21_6) + conv_s2u_18_19(data_rsci_idat[71:54]);
  assign MultLoop_acc_1385_nl = nl_MultLoop_acc_1385_nl[18:0];
  assign nl_MultLoop_acc_1325_nl =  -conv_s2s_13_14(data_rsci_idat[179:167]);
  assign MultLoop_acc_1325_nl = nl_MultLoop_acc_1325_nl[13:0];
  assign nl_MultLoop_acc_44_nl = conv_s2s_23_24({(~ (data_rsci_idat[179:162])) ,
      5'b00100}) + conv_s2s_20_24({(~ (data_rsci_idat[179:162])) , 2'b01}) + conv_s2s_19_24({(MultLoop_acc_1325_nl)
      , (~ (data_rsci_idat[166:162]))});
  assign MultLoop_acc_44_nl = nl_MultLoop_acc_44_nl[23:0];
  assign nl_MultLoop_acc_1085_nl = (readslicef_19_15_4((MultLoop_acc_1385_nl))) +
      conv_s2s_14_15(readslicef_24_14_10((MultLoop_acc_44_nl)));
  assign MultLoop_acc_1085_nl = nl_MultLoop_acc_1085_nl[14:0];
  assign nl_MultLoop_acc_34_nl = (MultLoop_acc_594_itm_18_2_1[16:6]) + 11'b00001010011;
  assign MultLoop_acc_34_nl = nl_MultLoop_acc_34_nl[10:0];
  assign nl_MultLoop_acc_1326_nl = conv_s2s_13_14(data_rsci_idat[35:23]) + 14'b00000000000001;
  assign MultLoop_acc_1326_nl = nl_MultLoop_acc_1326_nl[13:0];
  assign nl_MultLoop_acc_1069_nl = (~ (data_rsci_idat[35:18])) + conv_s2s_16_18({(MultLoop_acc_1326_nl)
      , (data_rsci_idat[22:21])});
  assign MultLoop_acc_1069_nl = nl_MultLoop_acc_1069_nl[17:0];
  assign nl_MultLoop_acc_298_nl = conv_s2u_18_21(MultLoop_acc_1069_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[35:18])) , 2'b01});
  assign MultLoop_acc_298_nl = nl_MultLoop_acc_298_nl[20:0];
  assign nl_MultLoop_22_MultLoop_acc_3_nl = conv_s2s_14_15({(MultLoop_acc_34_nl)
      , (MultLoop_acc_594_itm_18_2_1[5:3])}) + (readslicef_21_15_6((MultLoop_acc_298_nl)));
  assign MultLoop_22_MultLoop_acc_3_nl = nl_MultLoop_22_MultLoop_acc_3_nl[14:0];
  assign nl_MultLoop_acc_1072_nl = conv_s2s_18_19(data_rsci_idat[161:144]) + conv_s2s_13_19(data_rsci_idat[161:149]);
  assign MultLoop_acc_1072_nl = nl_MultLoop_acc_1072_nl[18:0];
  assign nl_MultLoop_acc_299_nl = conv_s2u_19_21(MultLoop_acc_1072_nl) + conv_s2u_20_21({(data_rsci_idat[161:144])
      , 2'b00});
  assign MultLoop_acc_299_nl = nl_MultLoop_acc_299_nl[20:0];
  assign nl_MultLoop_acc_1074_nl = ({(data_rsci_idat[89:72]) , 5'b00001}) + conv_s2s_19_23({Result_Result_conc_54_18_8
      , (~ (data_rsci_idat[79:72]))});
  assign MultLoop_acc_1074_nl = nl_MultLoop_acc_1074_nl[22:0];
  assign nl_MultLoop_acc_1322_nl = conv_s2u_15_18(readslicef_23_15_8((MultLoop_acc_1074_nl)))
      + (~ (data_rsci_idat[89:72]));
  assign MultLoop_acc_1322_nl = nl_MultLoop_acc_1322_nl[17:0];
  assign nl_MultLoop_acc_1091_nl = conv_s2s_17_18(MultLoop_acc_19_itm_19_3) + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_1324_nl)))
      + conv_s2s_15_18(MultLoop_acc_1085_nl) + conv_s2s_15_18(MultLoop_22_MultLoop_acc_3_nl)
      + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_299_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_1322_nl)));
  assign MultLoop_acc_1091_nl = nl_MultLoop_acc_1091_nl[17:0];
  assign nl_MultLoop_acc_1080_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_17_18({MultLoop_acc_1203_cse_1
      , (data_rsci_idat[45:38])});
  assign MultLoop_acc_1080_nl = nl_MultLoop_acc_1080_nl[17:0];
  assign nl_MultLoop_acc_1081_nl = conv_s2s_23_24({(~ (data_rsci_idat[53:36])) ,
      5'b00001}) + conv_s2s_18_24(MultLoop_acc_1080_nl);
  assign MultLoop_acc_1081_nl = nl_MultLoop_acc_1081_nl[23:0];
  assign nl_MultLoop_acc_37_nl = conv_s2u_24_26(MultLoop_acc_1081_nl) + ({(~ (data_rsci_idat[53:36]))
      , 8'b00100000});
  assign MultLoop_acc_37_nl = nl_MultLoop_acc_37_nl[25:0];
  assign nl_MultLoop_acc_1083_nl = ({(~ (data_rsci_idat[143:126])) , 5'b00000}) +
      conv_s2s_21_23(MultLoop_acc_623_cse_1);
  assign MultLoop_acc_1083_nl = nl_MultLoop_acc_1083_nl[22:0];
  assign nl_MultLoop_acc_1084_nl = conv_s2s_26_27({(~ (data_rsci_idat[143:126]))
      , 8'b00100000}) + conv_s2s_23_27(MultLoop_acc_1083_nl);
  assign MultLoop_acc_1084_nl = nl_MultLoop_acc_1084_nl[26:0];
  assign nl_MultLoop_acc_1328_nl = conv_s2u_19_20(readslicef_27_19_8((MultLoop_acc_1084_nl)))
      + ({(data_rsci_idat[143:126]) , 2'b01});
  assign MultLoop_acc_1328_nl = nl_MultLoop_acc_1328_nl[19:0];
  assign nl_MultLoop_acc_1090_nl = (readslicef_26_18_8((MultLoop_acc_37_nl))) + (readslicef_20_18_2((MultLoop_acc_1328_nl)));
  assign MultLoop_acc_1090_nl = nl_MultLoop_acc_1090_nl[17:0];
  assign nl_res_rsci_d_53_36  = (MultLoop_acc_1091_nl) + (MultLoop_acc_1090_nl);
  assign nl_Result_acc_37_nl = conv_s2s_24_25({(~ (data_rsci_idat[107:90])) , 6'b000100})
      + conv_s2s_20_25({(~ (data_rsci_idat[107:90])) , 2'b01}) + conv_s2s_19_25({Result_Result_conc_62_18_6
      , (~ (data_rsci_idat[95:90]))});
  assign Result_acc_37_nl = nl_Result_acc_37_nl[24:0];
  assign nl_Result_acc_146_nl = conv_s2s_22_23({(~ (data_rsci_idat[161:144])) , 4'b0100})
      + conv_s2s_21_23(MultLoop_acc_565_cse_1);
  assign Result_acc_146_nl = nl_Result_acc_146_nl[22:0];
  assign nl_Result_acc_40_nl = conv_s2s_23_24(Result_acc_146_nl) + ({(data_rsci_idat[161:144])
      , 6'b010000});
  assign Result_acc_40_nl = nl_Result_acc_40_nl[23:0];
  assign nl_MultLoop_acc_444_nl = conv_s2s_17_18(readslicef_25_17_8((Result_acc_37_nl)))
      + conv_s2s_17_18(readslicef_24_17_7((Result_acc_40_nl)));
  assign MultLoop_acc_444_nl = nl_MultLoop_acc_444_nl[17:0];
  assign nl_Result_acc_147_nl = (~ (data_rsci_idat[125:108])) + conv_s2s_13_18(data_rsci_idat[125:113]);
  assign Result_acc_147_nl = nl_Result_acc_147_nl[17:0];
  assign nl_Result_acc_44_nl = conv_s2u_18_20(Result_acc_147_nl) + ({(data_rsci_idat[125:108])
      , 2'b01});
  assign Result_acc_44_nl = nl_Result_acc_44_nl[19:0];
  assign nl_MultLoop_acc_447_nl = (MultLoop_acc_444_nl) + (readslicef_20_18_2((Result_acc_44_nl)));
  assign MultLoop_acc_447_nl = nl_MultLoop_acc_447_nl[17:0];
  assign nl_Result_acc_148_nl = ({(data_rsci_idat[143:126]) , 6'b000001}) + conv_s2s_18_24(~
      (data_rsci_idat[143:126]));
  assign Result_acc_148_nl = nl_Result_acc_148_nl[23:0];
  assign nl_Result_acc_217_nl = conv_s2u_16_19(readslicef_24_16_8((Result_acc_148_nl)))
      + conv_s2u_18_19(data_rsci_idat[143:126]);
  assign Result_acc_217_nl = nl_Result_acc_217_nl[18:0];
  assign nl_MultLoop_acc_1320_nl = conv_s2s_11_12(Result_acc_41_itm_20_8[12:2]) +
      12'b000001110011;
  assign MultLoop_acc_1320_nl = nl_MultLoop_acc_1320_nl[11:0];
  assign nl_Result_acc_35_nl = conv_s2u_16_18(data_rsci_idat[71:56]) - (data_rsci_idat[71:54]);
  assign Result_acc_35_nl = nl_Result_acc_35_nl[17:0];
  assign nl_Result_acc_42_nl = conv_s2u_15_19(data_rsci_idat[35:21]) + conv_s2u_18_19(data_rsci_idat[35:18]);
  assign Result_acc_42_nl = nl_Result_acc_42_nl[18:0];
  assign nl_MultLoop_acc_442_nl = conv_s2s_14_15({(MultLoop_acc_1320_nl) , (Result_acc_41_itm_20_8[1:0])})
      + conv_s2s_14_15(readslicef_18_14_4((Result_acc_35_nl))) + conv_s2s_13_15(readslicef_19_13_6((Result_acc_42_nl)));
  assign MultLoop_acc_442_nl = nl_MultLoop_acc_442_nl[14:0];
  assign nl_Result_acc_140_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_15_18({MultLoop_acc_1178_cse_1
      , (data_rsci_idat[41:40])});
  assign Result_acc_140_nl = nl_Result_acc_140_nl[17:0];
  assign nl_Result_acc_43_nl = conv_s2u_18_21(Result_acc_140_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[53:36])) , 2'b01});
  assign Result_acc_43_nl = nl_Result_acc_43_nl[20:0];
  assign nl_MultLoop_acc_443_nl = conv_s2s_15_17(MultLoop_acc_442_nl) + conv_s2s_16_17(readslicef_21_16_5((Result_acc_43_nl)));
  assign MultLoop_acc_443_nl = nl_MultLoop_acc_443_nl[16:0];
  assign nl_MultLoop_acc_446_nl = (readslicef_19_18_1((Result_acc_217_nl))) + conv_s2s_17_18(MultLoop_acc_443_nl);
  assign MultLoop_acc_446_nl = nl_MultLoop_acc_446_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_6_nl = conv_s2s_23_24({(~
      (data_rsci_idat[17:0])) , 5'b01000}) + conv_s2s_22_24(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_5_cse_1);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_6_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_6_nl[23:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_nl = conv_s2s_24_27(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_6_nl)
      + ({(data_rsci_idat[17:0]) , 9'b000100000});
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_nl[26:0];
  assign nl_Result_acc_220_nl =  -conv_s2s_11_12(data_rsci_idat[89:79]);
  assign Result_acc_220_nl = nl_Result_acc_220_nl[11:0];
  assign nl_Result_acc_142_nl = ({(data_rsci_idat[89:72]) , 2'b01}) + conv_s2s_19_20({(Result_acc_220_nl)
      , (~ (data_rsci_idat[78:72]))});
  assign Result_acc_142_nl = nl_Result_acc_142_nl[19:0];
  assign nl_Result_acc_221_nl = conv_s2u_13_18(readslicef_20_13_7((Result_acc_142_nl)))
      + (~ (data_rsci_idat[89:72]));
  assign Result_acc_221_nl = nl_Result_acc_221_nl[17:0];
  assign nl_res_rsci_d_521_504  = (MultLoop_acc_447_nl) + (MultLoop_acc_446_nl) +
      conv_s2s_17_18(readslicef_27_17_10((nnet_product_input_t_config2_weight_t_config2_accum_t_acc_nl)))
      + conv_s2s_17_18(readslicef_18_17_1((Result_acc_221_nl)));
  assign nl_MultLoop_acc_1044_nl = (~ (data_rsci_idat[125:108])) + conv_s2s_16_18({Result_acc_207_cse_1
      , (data_rsci_idat[114:111])});
  assign MultLoop_acc_1044_nl = nl_MultLoop_acc_1044_nl[17:0];
  assign nl_MultLoop_acc_1045_nl = conv_s2s_20_21({(~ (data_rsci_idat[125:108]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_1044_nl);
  assign MultLoop_acc_1045_nl = nl_MultLoop_acc_1045_nl[20:0];
  assign nl_MultLoop_acc_305_nl = conv_s2u_21_23(MultLoop_acc_1045_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[125:108])) , 4'b0100});
  assign MultLoop_acc_305_nl = nl_MultLoop_acc_305_nl[22:0];
  assign nl_MultLoop_acc_1317_nl =  -conv_s2s_13_14(data_rsci_idat[143:131]);
  assign MultLoop_acc_1317_nl = nl_MultLoop_acc_1317_nl[13:0];
  assign nl_MultLoop_acc_1047_nl = ({(data_rsci_idat[143:126]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_1317_nl)
      , (~ (data_rsci_idat[130:126]))});
  assign MultLoop_acc_1047_nl = nl_MultLoop_acc_1047_nl[20:0];
  assign nl_MultLoop_acc_53_nl = conv_s2s_21_23(MultLoop_acc_1047_nl) + ({(~ (data_rsci_idat[143:126]))
      , 5'b00000});
  assign MultLoop_acc_53_nl = nl_MultLoop_acc_53_nl[22:0];
  assign nl_MultLoop_acc_1063_nl = (MultLoop_acc_777_sdt_1[19:2]) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_305_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_53_nl)));
  assign MultLoop_acc_1063_nl = nl_MultLoop_acc_1063_nl[17:0];
  assign nl_MultLoop_acc_1412_nl = conv_s2u_18_20(MultLoop_acc_1395_itm_20_3_1) +
      ({(data_rsci_idat[53:36]) , 2'b01});
  assign MultLoop_acc_1412_nl = nl_MultLoop_acc_1412_nl[19:0];
  assign nl_MultLoop_acc_1319_nl = (MultLoop_acc_45_itm_22_9[13:3]) + 11'b00000001001;
  assign MultLoop_acc_1319_nl = nl_MultLoop_acc_1319_nl[10:0];
  assign nl_MultLoop_acc_1405_nl = conv_s2u_19_21(MultLoop_acc_1403_itm_20_2_1) +
      ({(data_rsci_idat[35:18]) , 3'b001});
  assign MultLoop_acc_1405_nl = nl_MultLoop_acc_1405_nl[20:0];
  assign nl_MultLoop_34_MultLoop_acc_3_nl = conv_s2s_16_17(readslicef_20_16_4((MultLoop_acc_1412_nl)))
      + conv_s2s_16_17(MultLoop_acc_302_itm_23_7[16:1]) + conv_s2s_14_17({(MultLoop_acc_1319_nl)
      , (MultLoop_acc_45_itm_22_9[2:0])}) + conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_1405_nl)));
  assign MultLoop_34_MultLoop_acc_3_nl = nl_MultLoop_34_MultLoop_acc_3_nl[16:0];
  assign nl_MultLoop_acc_1042_nl = (~ (data_rsci_idat[161:144])) + conv_s2s_14_18(data_rsci_idat[161:148]);
  assign MultLoop_acc_1042_nl = nl_MultLoop_acc_1042_nl[17:0];
  assign nl_MultLoop_acc_306_nl = conv_s2u_18_20(MultLoop_acc_1042_nl) + ({(data_rsci_idat[161:144])
      , 2'b01});
  assign MultLoop_acc_306_nl = nl_MultLoop_acc_306_nl[19:0];
  assign nl_MultLoop_acc_1065_nl = (MultLoop_acc_1063_nl) + conv_s2s_17_18(MultLoop_34_MultLoop_acc_3_nl)
      + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_306_nl)));
  assign MultLoop_acc_1065_nl = nl_MultLoop_acc_1065_nl[17:0];
  assign nl_MultLoop_acc_1058_nl = conv_s2s_22_23({(~ (data_rsci_idat[89:72])) ,
      4'b0100}) + conv_s2s_20_23({(~ (data_rsci_idat[89:72])) , 2'b01}) + conv_s2s_18_23(MultLoop_acc_1017_cse_1);
  assign MultLoop_acc_1058_nl = nl_MultLoop_acc_1058_nl[22:0];
  assign nl_MultLoop_acc_303_nl = conv_s2u_23_24(MultLoop_acc_1058_nl) + ({(data_rsci_idat[89:72])
      , 6'b010000});
  assign MultLoop_acc_303_nl = nl_MultLoop_acc_303_nl[23:0];
  assign nl_MultLoop_acc_1060_nl = conv_s2s_21_22({(data_rsci_idat[107:90]) , 3'b000})
      + conv_s2s_19_22(MultLoop_acc_405_cse_1);
  assign MultLoop_acc_1060_nl = nl_MultLoop_acc_1060_nl[21:0];
  assign nl_MultLoop_acc_304_nl = conv_s2u_22_24(MultLoop_acc_1060_nl) + conv_s2u_23_24({(data_rsci_idat[107:90])
      , 5'b00000});
  assign MultLoop_acc_304_nl = nl_MultLoop_acc_304_nl[23:0];
  assign nl_MultLoop_acc_1064_nl = (readslicef_24_18_6((MultLoop_acc_303_nl))) +
      (readslicef_24_18_6((MultLoop_acc_304_nl)));
  assign MultLoop_acc_1064_nl = nl_MultLoop_acc_1064_nl[17:0];
  assign nl_res_rsci_d_71_54  = (MultLoop_acc_1065_nl) + (MultLoop_acc_1064_nl);
  assign nl_Result_acc_162_nl = conv_s2s_23_24({(~ (data_rsci_idat[71:54])) , 5'b01000})
      + conv_s2s_22_24(MultLoop_acc_473_cse_1);
  assign Result_acc_162_nl = nl_Result_acc_162_nl[23:0];
  assign nl_Result_acc_23_nl = conv_s2s_24_25(Result_acc_162_nl) + ({(data_rsci_idat[71:54])
      , 7'b0100000});
  assign Result_acc_23_nl = nl_Result_acc_23_nl[24:0];
  assign nl_Result_acc_28_nl = conv_s2s_26_27({(~ (data_rsci_idat[161:144])) , 8'b00100000})
      + conv_s2s_23_27({(~ (data_rsci_idat[161:144])) , 5'b00100}) + conv_s2s_21_27(MultLoop_acc_763_cse_1);
  assign Result_acc_28_nl = nl_Result_acc_28_nl[26:0];
  assign nl_MultLoop_acc_455_nl = (readslicef_25_18_7((Result_acc_23_nl))) + (readslicef_27_18_9((Result_acc_28_nl)));
  assign MultLoop_acc_455_nl = nl_MultLoop_acc_455_nl[17:0];
  assign nl_Result_acc_155_nl = ({(data_rsci_idat[53:36]) , 4'b0001}) + conv_s2s_18_22(~
      (data_rsci_idat[53:36]));
  assign Result_acc_155_nl = nl_Result_acc_155_nl[21:0];
  assign nl_Result_acc_212_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_16_18(readslicef_22_16_6((Result_acc_155_nl)));
  assign Result_acc_212_nl = nl_Result_acc_212_nl[17:0];
  assign nl_Result_acc_213_nl = conv_s2u_18_20(Result_acc_212_nl) + ({(data_rsci_idat[53:36])
      , 2'b01});
  assign Result_acc_213_nl = nl_Result_acc_213_nl[19:0];
  assign nl_Result_acc_25_nl = conv_s2u_15_18(data_rsci_idat[107:93]) - (data_rsci_idat[107:90]);
  assign Result_acc_25_nl = nl_Result_acc_25_nl[17:0];
  assign nl_Result_acc_24_nl = conv_s2s_24_25({(~ (data_rsci_idat[89:72])) , 6'b010000})
      + conv_s2s_22_25({(~ (data_rsci_idat[89:72])) , 4'b0100}) + conv_s2s_20_25({(~
      (data_rsci_idat[89:72])) , 2'b01}) + conv_s2s_19_25({Result_Result_conc_56_18_6
      , (~ (data_rsci_idat[77:72]))});
  assign Result_acc_24_nl = nl_Result_acc_24_nl[24:0];
  assign nl_MultLoop_acc_454_nl = conv_s2s_17_18(readslicef_20_17_3((Result_acc_213_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((Result_acc_25_nl))) + conv_s2s_15_18(readslicef_25_15_10((Result_acc_24_nl)));
  assign MultLoop_acc_454_nl = nl_MultLoop_acc_454_nl[17:0];
  assign nl_MultLoop_acc_457_nl = (MultLoop_acc_455_nl) + (MultLoop_acc_454_nl);
  assign MultLoop_acc_457_nl = nl_MultLoop_acc_457_nl[17:0];
  assign nl_Result_acc_158_nl = conv_s2s_18_19(data_rsci_idat[143:126]) + conv_s2s_14_19({Result_acc_202_cse_1
      , (data_rsci_idat[134:131])});
  assign Result_acc_158_nl = nl_Result_acc_158_nl[18:0];
  assign nl_Result_acc_27_nl = conv_s2u_19_22(Result_acc_158_nl) + ({(~ (data_rsci_idat[143:126]))
      , 4'b0000});
  assign Result_acc_27_nl = nl_Result_acc_27_nl[21:0];
  assign nl_Result_acc_154_nl = conv_s2s_21_22({(~ (data_rsci_idat[179:162])) , 3'b001})
      + conv_s2s_18_22(Result_acc_195_cse_1);
  assign Result_acc_154_nl = nl_Result_acc_154_nl[21:0];
  assign nl_Result_acc_31_nl = conv_s2u_22_23(Result_acc_154_nl) + ({(data_rsci_idat[179:162])
      , 5'b01000});
  assign Result_acc_31_nl = nl_Result_acc_31_nl[22:0];
  assign nl_Result_acc_215_nl =  -conv_s2s_16_17(data_rsci_idat[35:20]);
  assign Result_acc_215_nl = nl_Result_acc_215_nl[16:0];
  assign nl_Result_acc_21_nl = conv_s2s_19_21({(Result_acc_215_nl) , (~ (data_rsci_idat[19:18]))})
      + conv_s2s_20_21({(~ (data_rsci_idat[35:18])) , 2'b01});
  assign Result_acc_21_nl = nl_Result_acc_21_nl[20:0];
  assign nl_MultLoop_acc_449_nl = (readslicef_21_11_10((Result_acc_21_nl))) + 11'b00001101111;
  assign MultLoop_acc_449_nl = nl_MultLoop_acc_449_nl[10:0];
  assign nl_MultLoop_acc_450_nl = (MultLoop_acc_650_cse_1[18:7]) + conv_s2s_11_12(MultLoop_acc_449_nl);
  assign MultLoop_acc_450_nl = nl_MultLoop_acc_450_nl[11:0];
  assign nl_MultLoop_acc_453_nl = conv_s2s_17_18(readslicef_22_17_5((Result_acc_27_nl)))
      + conv_s2s_15_18(readslicef_23_15_8((Result_acc_31_nl))) + conv_s2s_12_18(MultLoop_acc_450_nl);
  assign MultLoop_acc_453_nl = nl_MultLoop_acc_453_nl[17:0];
  assign nl_Result_acc_160_nl = (~ (data_rsci_idat[17:0])) + conv_s2s_17_18({MultLoop_acc_1151_cse_1
      , (data_rsci_idat[7:2])});
  assign Result_acc_160_nl = nl_Result_acc_160_nl[17:0];
  assign nl_Result_acc_32_nl = conv_s2u_18_25(Result_acc_160_nl) + conv_s2u_24_25({(~
      (data_rsci_idat[17:0])) , 6'b000001});
  assign Result_acc_32_nl = nl_Result_acc_32_nl[24:0];
  assign nl_MultLoop_acc_456_nl = (MultLoop_acc_453_nl) + (readslicef_25_18_7((Result_acc_32_nl)));
  assign MultLoop_acc_456_nl = nl_MultLoop_acc_456_nl[17:0];
  assign nl_res_rsci_d_503_486  = (MultLoop_acc_457_nl) + (MultLoop_acc_456_nl);
  assign nl_MultLoop_acc_1384_nl = ({(data_rsci_idat[125:108]) , 4'b0001}) + conv_s2u_19_22(MultLoop_acc_808_itm_20_2_1);
  assign MultLoop_acc_1384_nl = nl_MultLoop_acc_1384_nl[21:0];
  assign nl_MultLoop_acc_1313_nl = conv_s2u_16_19(readslicef_22_16_6((MultLoop_acc_1384_nl)))
      + conv_s2u_18_19(data_rsci_idat[125:108]);
  assign MultLoop_acc_1313_nl = nl_MultLoop_acc_1313_nl[18:0];
  assign nl_MultLoop_acc_1030_nl = ({(data_rsci_idat[53:36]) , 6'b010000}) + conv_s2s_22_24({(~
      (data_rsci_idat[53:36])) , 4'b0100}) + conv_s2s_21_24(MultLoop_acc_789_cse_1);
  assign MultLoop_acc_1030_nl = nl_MultLoop_acc_1030_nl[23:0];
  assign nl_MultLoop_acc_1315_nl = conv_s2u_16_18(readslicef_24_16_8((MultLoop_acc_1030_nl)))
      + (~ (data_rsci_idat[53:36]));
  assign MultLoop_acc_1315_nl = nl_MultLoop_acc_1315_nl[17:0];
  assign nl_MultLoop_acc_57_nl = (MultLoop_acc_56_itm_17_1[16:1]) + 16'b0000000011010001;
  assign MultLoop_acc_57_nl = nl_MultLoop_acc_57_nl[15:0];
  assign nl_MultLoop_acc_1016_nl = (~ (data_rsci_idat[143:126])) + conv_s2s_14_18(data_rsci_idat[143:130]);
  assign MultLoop_acc_1016_nl = nl_MultLoop_acc_1016_nl[17:0];
  assign nl_MultLoop_acc_310_nl = conv_s2u_18_21(MultLoop_acc_1016_nl) + ({(data_rsci_idat[143:126])
      , 3'b001});
  assign MultLoop_acc_310_nl = nl_MultLoop_acc_310_nl[20:0];
  assign nl_MultLoop_acc_1040_nl = conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_1313_nl)))
      + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_1315_nl))) + conv_s2s_17_18({(MultLoop_acc_57_nl)
      , (MultLoop_acc_56_itm_17_1[0])}) + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_310_nl)));
  assign MultLoop_acc_1040_nl = nl_MultLoop_acc_1040_nl[17:0];
  assign nl_MultLoop_acc_1309_nl = conv_s2s_11_12(data_rsci_idat[107:97]) + 12'b000000000001;
  assign MultLoop_acc_1309_nl = nl_MultLoop_acc_1309_nl[11:0];
  assign nl_MultLoop_acc_1032_nl = (~ (data_rsci_idat[107:90])) + conv_s2s_17_18({(MultLoop_acc_1309_nl)
      , (data_rsci_idat[96:92])});
  assign MultLoop_acc_1032_nl = nl_MultLoop_acc_1032_nl[17:0];
  assign nl_MultLoop_acc_1033_nl = conv_s2s_21_22({(~ (data_rsci_idat[107:90])) ,
      3'b001}) + conv_s2s_18_22(MultLoop_acc_1032_nl);
  assign MultLoop_acc_1033_nl = nl_MultLoop_acc_1033_nl[21:0];
  assign nl_MultLoop_acc_309_nl = conv_s2u_22_24(MultLoop_acc_1033_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[107:90])) , 5'b01000});
  assign MultLoop_acc_309_nl = nl_MultLoop_acc_309_nl[23:0];
  assign nl_MultLoop_acc_308_nl = conv_s2u_18_21(MultLoop_acc_1017_cse_1) + ({(data_rsci_idat[89:72])
      , 3'b001});
  assign MultLoop_acc_308_nl = nl_MultLoop_acc_308_nl[20:0];
  assign nl_MultLoop_acc_1310_nl = conv_s2s_14_15(data_rsci_idat[71:58]) + 15'b000000000000001;
  assign MultLoop_acc_1310_nl = nl_MultLoop_acc_1310_nl[14:0];
  assign nl_MultLoop_acc_1019_nl = conv_s2s_18_19(data_rsci_idat[71:54]) + conv_s2s_17_19({(MultLoop_acc_1310_nl)
      , (data_rsci_idat[57:56])});
  assign MultLoop_acc_1019_nl = nl_MultLoop_acc_1019_nl[18:0];
  assign nl_MultLoop_acc_60_nl = conv_s2u_19_20(MultLoop_acc_1019_nl) + ({(~ (data_rsci_idat[71:54]))
      , 2'b00});
  assign MultLoop_acc_60_nl = nl_MultLoop_acc_60_nl[19:0];
  assign nl_MultLoop_acc_1035_nl = conv_s2s_16_17(readslicef_21_16_5((MultLoop_acc_308_nl)))
      + conv_s2s_16_17(readslicef_20_16_4((MultLoop_acc_60_nl)));
  assign MultLoop_acc_1035_nl = nl_MultLoop_acc_1035_nl[16:0];
  assign nl_MultLoop_acc_1039_nl = (readslicef_24_18_6((MultLoop_acc_309_nl))) +
      conv_s2s_17_18(MultLoop_acc_1035_nl);
  assign MultLoop_acc_1039_nl = nl_MultLoop_acc_1039_nl[17:0];
  assign nl_MultLoop_acc_1023_nl = ({(~ (data_rsci_idat[179:162])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_777_sdt_1);
  assign MultLoop_acc_1023_nl = nl_MultLoop_acc_1023_nl[21:0];
  assign nl_MultLoop_acc_1024_nl = ({(data_rsci_idat[179:162]) , 6'b010000}) + conv_s2s_22_24(MultLoop_acc_1023_nl);
  assign MultLoop_acc_1024_nl = nl_MultLoop_acc_1024_nl[23:0];
  assign nl_MultLoop_acc_1312_nl = conv_s2u_16_19(readslicef_24_16_8((MultLoop_acc_1024_nl)))
      + conv_s2u_18_19(data_rsci_idat[179:162]);
  assign MultLoop_acc_1312_nl = nl_MultLoop_acc_1312_nl[18:0];
  assign nl_MultLoop_acc_1021_nl = conv_s2s_20_21({(~ (data_rsci_idat[35:18])) ,
      2'b01}) + conv_s2s_18_21(MultLoop_acc_557_cse_1);
  assign MultLoop_acc_1021_nl = nl_MultLoop_acc_1021_nl[20:0];
  assign nl_MultLoop_acc_307_nl = conv_s2u_21_22(MultLoop_acc_1021_nl) + ({(data_rsci_idat[35:18])
      , 4'b0100});
  assign MultLoop_acc_307_nl = nl_MultLoop_acc_307_nl[21:0];
  assign nl_MultLoop_acc_65_nl = conv_s2s_24_25({(~ (data_rsci_idat[161:144])) ,
      6'b001000}) + conv_s2s_21_25({(~ (data_rsci_idat[161:144])) , 3'b001}) + conv_s2s_19_25({MultLoop_MultLoop_conc_212_18_6
      , (~ (data_rsci_idat[149:144]))});
  assign MultLoop_acc_65_nl = nl_MultLoop_acc_65_nl[24:0];
  assign nl_res_rsci_d_89_72  = (MultLoop_acc_1040_nl) + (MultLoop_acc_1039_nl) +
      conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_1312_nl))) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_307_nl)))
      + conv_s2s_15_18(readslicef_25_15_10((MultLoop_acc_65_nl)));
  assign nl_Result_acc_252_nl = conv_s2u_18_21(MultLoop_acc_1395_itm_20_3_1) + ({(data_rsci_idat[53:36])
      , 3'b001});
  assign Result_acc_252_nl = nl_Result_acc_252_nl[20:0];
  assign nl_Result_acc_170_nl = conv_s2s_18_19(data_rsci_idat[89:72]) + conv_s2s_15_19({MultLoop_acc_1150_cse_1
      , (data_rsci_idat[79:76])});
  assign Result_acc_170_nl = nl_Result_acc_170_nl[18:0];
  assign nl_Result_acc_9_nl = conv_s2u_19_22(Result_acc_170_nl) + ({(~ (data_rsci_idat[89:72]))
      , 4'b0000});
  assign Result_acc_9_nl = nl_Result_acc_9_nl[21:0];
  assign nl_MultLoop_acc_462_nl = conv_s2s_17_18(readslicef_21_17_4((Result_acc_252_nl)))
      + conv_s2s_16_18(readslicef_22_16_6((Result_acc_9_nl)));
  assign MultLoop_acc_462_nl = nl_MultLoop_acc_462_nl[17:0];
  assign nl_Result_acc_253_nl = conv_s2u_19_23(MultLoop_acc_1403_itm_20_2_1) + ({(data_rsci_idat[35:18])
      , 5'b00001});
  assign Result_acc_253_nl = nl_Result_acc_253_nl[22:0];
  assign nl_MultLoop_acc_465_nl = (MultLoop_acc_462_nl) + (readslicef_23_18_5((Result_acc_253_nl)));
  assign MultLoop_acc_465_nl = nl_MultLoop_acc_465_nl[17:0];
  assign nl_Result_acc_203_nl =  -conv_s2s_9_10(data_rsci_idat[161:153]);
  assign Result_acc_203_nl = nl_Result_acc_203_nl[9:0];
  assign nl_Result_acc_185_nl = ({(data_rsci_idat[161:144]) , 2'b01}) + conv_s2s_19_20({(Result_acc_203_nl)
      , (~ (data_rsci_idat[152:144]))});
  assign Result_acc_185_nl = nl_Result_acc_185_nl[19:0];
  assign nl_Result_acc_186_nl = conv_s2s_22_23({(data_rsci_idat[161:144]) , 4'b0000})
      + conv_s2s_20_23(Result_acc_185_nl);
  assign Result_acc_186_nl = nl_Result_acc_186_nl[22:0];
  assign nl_Result_acc_204_nl = (~ (data_rsci_idat[161:144])) + conv_s2s_16_18(readslicef_23_16_7((Result_acc_186_nl)));
  assign Result_acc_204_nl = nl_Result_acc_204_nl[17:0];
  assign nl_Result_acc_205_nl = conv_s2u_18_21(Result_acc_204_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[161:144])) , 2'b01});
  assign Result_acc_205_nl = nl_Result_acc_205_nl[20:0];
  assign nl_Result_acc_206_nl =  -conv_s2s_14_15(data_rsci_idat[107:94]);
  assign Result_acc_206_nl = nl_Result_acc_206_nl[14:0];
  assign nl_Result_acc_10_nl = conv_s2s_19_23({(Result_acc_206_nl) , (~ (data_rsci_idat[93:90]))})
      + conv_s2s_22_23({(~ (data_rsci_idat[107:90])) , 4'b0001});
  assign Result_acc_10_nl = nl_Result_acc_10_nl[22:0];
  assign nl_Result_acc_174_nl = conv_s2s_21_22({(data_rsci_idat[125:108]) , 3'b000})
      + conv_s2s_18_22(data_rsci_idat[125:108]) + conv_s2s_17_22({Result_acc_207_cse_1
      , (data_rsci_idat[114:110])});
  assign Result_acc_174_nl = nl_Result_acc_174_nl[21:0];
  assign nl_Result_acc_11_nl = conv_s2u_22_23(Result_acc_174_nl) + ({(~ (data_rsci_idat[125:108]))
      , 5'b00000});
  assign Result_acc_11_nl = nl_Result_acc_11_nl[22:0];
  assign nl_MultLoop_acc_461_nl = conv_s2s_16_17(readslicef_23_16_7((Result_acc_10_nl)))
      + conv_s2s_16_17(readslicef_23_16_7((Result_acc_11_nl)));
  assign MultLoop_acc_461_nl = nl_MultLoop_acc_461_nl[16:0];
  assign nl_MultLoop_acc_464_nl = (readslicef_21_18_3((Result_acc_205_nl))) + conv_s2s_17_18(MultLoop_acc_461_nl);
  assign MultLoop_acc_464_nl = nl_MultLoop_acc_464_nl[17:0];
  assign nl_Result_acc_179_nl = conv_s2s_22_23({(~ (data_rsci_idat[17:0])) , 4'b0100})
      + conv_s2s_20_23({(~ (data_rsci_idat[17:0])) , 2'b01}) + conv_s2s_18_23(MultLoop_acc_412_cse_1);
  assign Result_acc_179_nl = nl_Result_acc_179_nl[22:0];
  assign nl_Result_acc_17_nl = conv_s2u_23_24(Result_acc_179_nl) + ({(data_rsci_idat[17:0])
      , 6'b010000});
  assign Result_acc_17_nl = nl_Result_acc_17_nl[23:0];
  assign nl_Result_acc_176_nl = conv_s2s_20_21({(data_rsci_idat[143:126]) , 2'b00})
      + conv_s2s_19_21(Result_acc_175_cse);
  assign Result_acc_176_nl = nl_Result_acc_176_nl[20:0];
  assign nl_Result_acc_16_nl = conv_s2u_21_23(Result_acc_176_nl) + conv_s2u_22_23({(data_rsci_idat[143:126])
      , 4'b0000});
  assign Result_acc_16_nl = nl_Result_acc_16_nl[22:0];
  assign nl_Result_acc_208_nl =  -conv_s2s_13_14(data_rsci_idat[71:59]);
  assign Result_acc_208_nl = nl_Result_acc_208_nl[13:0];
  assign nl_Result_acc_167_nl = ({(data_rsci_idat[71:54]) , 2'b01}) + conv_s2s_19_20({(Result_acc_208_nl)
      , (~ (data_rsci_idat[58:54]))});
  assign Result_acc_167_nl = nl_Result_acc_167_nl[19:0];
  assign nl_Result_acc_8_nl = conv_s2s_20_23(Result_acc_167_nl) + ({(~ (data_rsci_idat[71:54]))
      , 5'b00000});
  assign Result_acc_8_nl = nl_Result_acc_8_nl[22:0];
  assign nl_MultLoop_acc_458_nl = conv_s2s_13_14(readslicef_23_13_10((Result_acc_8_nl)))
      + 14'b00000110111011;
  assign MultLoop_acc_458_nl = nl_MultLoop_acc_458_nl[13:0];
  assign nl_Result_acc_168_nl = (~ (data_rsci_idat[179:162])) + conv_s2s_14_18(data_rsci_idat[179:166]);
  assign Result_acc_168_nl = nl_Result_acc_168_nl[17:0];
  assign nl_Result_acc_15_nl = conv_s2u_18_20(Result_acc_168_nl) + ({(data_rsci_idat[179:162])
      , 2'b01});
  assign Result_acc_15_nl = nl_Result_acc_15_nl[19:0];
  assign nl_res_rsci_d_485_468  = (MultLoop_acc_465_nl) + (MultLoop_acc_464_nl) +
      conv_s2s_17_18(readslicef_24_17_7((Result_acc_17_nl))) + conv_s2s_16_18(readslicef_23_16_7((Result_acc_16_nl)))
      + conv_s2s_14_18(MultLoop_acc_458_nl) + conv_s2s_14_18(readslicef_20_14_6((Result_acc_15_nl)));
  assign nl_MultLoop_acc_1005_nl = conv_s2s_22_23({(~ (data_rsci_idat[71:54])) ,
      4'b0001}) + conv_s2s_18_23(MultLoop_acc_410_cse_1);
  assign MultLoop_acc_1005_nl = nl_MultLoop_acc_1005_nl[22:0];
  assign nl_MultLoop_acc_311_nl = conv_s2u_23_24(MultLoop_acc_1005_nl) + ({(data_rsci_idat[71:54])
      , 6'b010000});
  assign MultLoop_acc_311_nl = nl_MultLoop_acc_311_nl[23:0];
  assign nl_MultLoop_acc_1394_nl = conv_s2u_18_22(MultLoop_asn_361) + ({(data_rsci_idat[179:162])
      , 4'b0001});
  assign MultLoop_acc_1394_nl = nl_MultLoop_acc_1394_nl[21:0];
  assign nl_MultLoop_acc_75_nl = conv_s2u_13_18(data_rsci_idat[161:149]) - (data_rsci_idat[161:144]);
  assign MultLoop_acc_75_nl = nl_MultLoop_acc_75_nl[17:0];
  assign nl_MultLoop_acc_1383_nl = conv_s2u_19_20(MultLoop_acc_839_cse_1[21:3]) +
      ({(data_rsci_idat[35:18]) , 2'b01});
  assign MultLoop_acc_1383_nl = nl_MultLoop_acc_1383_nl[19:0];
  assign nl_MultLoop_acc_1006_nl = (readslicef_20_14_6((MultLoop_acc_1383_nl))) +
      conv_s2s_11_14(MultLoop_acc_405_cse_1[18:8]);
  assign MultLoop_acc_1006_nl = nl_MultLoop_acc_1006_nl[13:0];
  assign nl_MultLoop_acc_1302_nl =  -conv_s2s_13_14(data_rsci_idat[125:113]);
  assign MultLoop_acc_1302_nl = nl_MultLoop_acc_1302_nl[13:0];
  assign nl_MultLoop_acc_73_nl = conv_s2s_23_24({(~ (data_rsci_idat[125:108])) ,
      5'b00100}) + conv_s2s_20_24({(~ (data_rsci_idat[125:108])) , 2'b01}) + conv_s2s_19_24({(MultLoop_acc_1302_nl)
      , (~ (data_rsci_idat[112:108]))});
  assign MultLoop_acc_73_nl = nl_MultLoop_acc_73_nl[23:0];
  assign nl_MultLoop_acc_1009_nl = conv_s2s_16_17(readslicef_22_16_6((MultLoop_acc_1394_nl)))
      + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_75_nl))) + conv_s2s_14_17(MultLoop_acc_1006_nl)
      + conv_s2s_14_17(readslicef_24_14_10((MultLoop_acc_73_nl)));
  assign MultLoop_acc_1009_nl = nl_MultLoop_acc_1009_nl[16:0];
  assign nl_MultLoop_acc_1011_nl = (readslicef_24_18_6((MultLoop_acc_311_nl))) +
      conv_s2s_17_18(MultLoop_acc_1009_nl);
  assign MultLoop_acc_1011_nl = nl_MultLoop_acc_1011_nl[17:0];
  assign nl_MultLoop_acc_1304_nl = conv_s2u_18_19(data_rsci_idat[89:72]) + conv_s2u_14_19(MultLoop_acc_1399_itm_20_5[15:2]);
  assign MultLoop_acc_1304_nl = nl_MultLoop_acc_1304_nl[18:0];
  assign nl_MultLoop_acc_1305_nl = conv_s2u_17_18(readslicef_19_17_2((MultLoop_acc_1304_nl)))
      + (~ (data_rsci_idat[89:72]));
  assign MultLoop_acc_1305_nl = nl_MultLoop_acc_1305_nl[17:0];
  assign nl_MultLoop_acc_1013_nl = (MultLoop_acc_1011_nl) + conv_s2s_17_18(MultLoop_acc_74_itm_17_1)
      + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_1305_nl)));
  assign MultLoop_acc_1013_nl = nl_MultLoop_acc_1013_nl[17:0];
  assign nl_MultLoop_acc_1000_nl = ({(data_rsci_idat[17:0]) , 4'b0100}) + conv_s2s_21_22(MultLoop_acc_744_cse_1);
  assign MultLoop_acc_1000_nl = nl_MultLoop_acc_1000_nl[21:0];
  assign nl_MultLoop_acc_1001_nl = conv_s2s_24_25({(data_rsci_idat[17:0]) , 6'b000000})
      + conv_s2s_22_25(MultLoop_acc_1000_nl);
  assign MultLoop_acc_1001_nl = nl_MultLoop_acc_1001_nl[24:0];
  assign nl_MultLoop_acc_1306_nl = conv_s2u_17_19(readslicef_25_17_8((MultLoop_acc_1001_nl)))
      + conv_s2u_18_19(data_rsci_idat[17:0]);
  assign MultLoop_acc_1306_nl = nl_MultLoop_acc_1306_nl[18:0];
  assign nl_MultLoop_acc_1307_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_14_18(MultLoop_acc_596_itm_20_5[15:2]);
  assign MultLoop_acc_1307_nl = nl_MultLoop_acc_1307_nl[17:0];
  assign nl_MultLoop_acc_1308_nl = conv_s2u_18_20(MultLoop_acc_1307_nl) + ({(data_rsci_idat[53:36])
      , 2'b01});
  assign MultLoop_acc_1308_nl = nl_MultLoop_acc_1308_nl[19:0];
  assign nl_MultLoop_acc_1012_nl = (readslicef_19_18_1((MultLoop_acc_1306_nl))) +
      (readslicef_20_18_2((MultLoop_acc_1308_nl)));
  assign MultLoop_acc_1012_nl = nl_MultLoop_acc_1012_nl[17:0];
  assign nl_res_rsci_d_107_90  = (MultLoop_acc_1013_nl) + (MultLoop_acc_1012_nl);
  assign nl_Result_acc_250_nl = conv_s2u_18_19(data_rsci_idat[161:144]) + conv_s2u_16_19(MultLoop_acc_714_itm_19_4);
  assign Result_acc_250_nl = nl_Result_acc_250_nl[18:0];
  assign nl_Result_acc_199_nl = conv_s2u_15_18(readslicef_19_15_4((Result_acc_250_nl)))
      + (~ (data_rsci_idat[161:144]));
  assign Result_acc_199_nl = nl_Result_acc_199_nl[17:0];
  assign nl_MultLoop_acc_1381_nl = conv_s2u_19_20(MultLoop_acc_473_cse_1[21:3]) +
      ({(data_rsci_idat[71:54]) , 2'b01});
  assign MultLoop_acc_1381_nl = nl_MultLoop_acc_1381_nl[19:0];
  assign nl_MultLoop_acc_477_nl = conv_s2s_17_18(readslicef_18_17_1((Result_acc_199_nl)))
      + conv_s2s_17_18(readslicef_20_17_3((MultLoop_acc_1381_nl)));
  assign MultLoop_acc_477_nl = nl_MultLoop_acc_477_nl[17:0];
  assign nl_MultLoop_acc_1382_nl = conv_s2u_18_19(data_rsci_idat[53:36]) + conv_s2u_16_19(MultLoop_acc_733_cse_1[19:4]);
  assign MultLoop_acc_1382_nl = nl_MultLoop_acc_1382_nl[18:0];
  assign nl_MultLoop_acc_1298_nl = conv_s2u_15_19(readslicef_19_15_4((MultLoop_acc_1382_nl)))
      + conv_s2u_18_19(data_rsci_idat[53:36]);
  assign MultLoop_acc_1298_nl = nl_MultLoop_acc_1298_nl[18:0];
  assign nl_MultLoop_acc_481_nl = (MultLoop_acc_477_nl) + (readslicef_19_18_1((MultLoop_acc_1298_nl)));
  assign MultLoop_acc_481_nl = nl_MultLoop_acc_481_nl[17:0];
  assign nl_Result_acc_194_nl = ({(data_rsci_idat[125:108]) , 6'b000001}) + conv_s2s_18_24(~
      (data_rsci_idat[125:108]));
  assign Result_acc_194_nl = nl_Result_acc_194_nl[23:0];
  assign nl_Result_acc_nl = conv_s2u_16_19(readslicef_24_16_8((Result_acc_194_nl)))
      + conv_s2u_18_19(data_rsci_idat[125:108]);
  assign Result_acc_nl = nl_Result_acc_nl[18:0];
  assign nl_Result_acc_196_nl = ({(data_rsci_idat[179:162]) , 4'b0001}) + conv_s2s_18_22(Result_acc_195_cse_1);
  assign Result_acc_196_nl = nl_Result_acc_196_nl[21:0];
  assign nl_Result_acc_200_nl = (~ (data_rsci_idat[179:162])) + conv_s2s_16_18(readslicef_22_16_6((Result_acc_196_nl)));
  assign Result_acc_200_nl = nl_Result_acc_200_nl[17:0];
  assign nl_Result_acc_201_nl = conv_s2u_18_20(Result_acc_200_nl) + ({(data_rsci_idat[179:162])
      , 2'b01});
  assign Result_acc_201_nl = nl_Result_acc_201_nl[19:0];
  assign nl_MultLoop_acc_480_nl = (readslicef_19_18_1((Result_acc_nl))) + (readslicef_20_18_2((Result_acc_201_nl)));
  assign MultLoop_acc_480_nl = nl_MultLoop_acc_480_nl[17:0];
  assign nl_MultLoop_acc_483_nl = (MultLoop_acc_481_nl) + (MultLoop_acc_480_nl);
  assign MultLoop_acc_483_nl = nl_MultLoop_acc_483_nl[17:0];
  assign nl_MultLoop_acc_469_nl = (~ (data_rsci_idat[89:72])) + conv_s2s_17_18({MultLoop_acc_1150_cse_1
      , (data_rsci_idat[79:74])});
  assign MultLoop_acc_469_nl = nl_MultLoop_acc_469_nl[17:0];
  assign nl_MultLoop_acc_470_nl = ({(data_rsci_idat[89:72]) , 4'b0001}) + conv_s2s_18_22(MultLoop_acc_469_nl);
  assign MultLoop_acc_470_nl = nl_MultLoop_acc_470_nl[21:0];
  assign nl_MultLoop_acc_1301_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_470_nl)))
      + (~ (data_rsci_idat[89:72]));
  assign MultLoop_acc_1301_nl = nl_MultLoop_acc_1301_nl[17:0];
  assign nl_MultLoop_acc_467_nl = ({(data_rsci_idat[35:18]) , 4'b0001}) + conv_s2s_18_22(~
      (data_rsci_idat[35:18]));
  assign MultLoop_acc_467_nl = nl_MultLoop_acc_467_nl[21:0];
  assign nl_MultLoop_acc_1299_nl = conv_s2u_15_19(readslicef_22_15_7((MultLoop_acc_467_nl)))
      + conv_s2u_18_19(data_rsci_idat[35:18]);
  assign MultLoop_acc_1299_nl = nl_MultLoop_acc_1299_nl[18:0];
  assign nl_MultLoop_acc_278_nl = (MultLoop_acc_279_itm_20_6[14:1]) + 14'b11111111111101;
  assign MultLoop_acc_278_nl = nl_MultLoop_acc_278_nl[13:0];
  assign nl_MultLoop_acc_472_nl = conv_s2s_24_25({(~ (data_rsci_idat[107:90])) ,
      6'b000100}) + conv_s2s_20_25({(~ (data_rsci_idat[107:90])) , 2'b01}) + conv_s2s_18_25(~
      (data_rsci_idat[107:90]));
  assign MultLoop_acc_472_nl = nl_MultLoop_acc_472_nl[24:0];
  assign nl_MultLoop_acc_284_nl = conv_s2s_25_26(MultLoop_acc_472_nl) + ({(data_rsci_idat[107:90])
      , 8'b01000000});
  assign MultLoop_acc_284_nl = nl_MultLoop_acc_284_nl[25:0];
  assign nl_Result_acc_189_nl = (~ (data_rsci_idat[143:126])) + conv_s2s_15_18({Result_acc_202_cse_1
      , (data_rsci_idat[134:130])});
  assign Result_acc_189_nl = nl_Result_acc_189_nl[17:0];
  assign nl_Result_acc_190_nl = ({(data_rsci_idat[143:126]) , 3'b001}) + conv_s2s_18_21(Result_acc_189_nl);
  assign Result_acc_190_nl = nl_Result_acc_190_nl[20:0];
  assign nl_Result_acc_2_nl = conv_s2u_21_23(Result_acc_190_nl) + ({(~ (data_rsci_idat[143:126]))
      , 5'b00000});
  assign Result_acc_2_nl = nl_Result_acc_2_nl[22:0];
  assign nl_res_rsci_d_467_450  = (MultLoop_acc_483_nl) + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_1301_nl)))
      + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_1299_nl))) + conv_s2s_15_18({(MultLoop_acc_278_nl)
      , (MultLoop_acc_279_itm_20_6[0])}) + conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_284_nl)))
      + conv_s2s_17_18(readslicef_23_17_6((Result_acc_2_nl)));
  assign nl_MultLoop_acc_1380_nl = conv_s2u_18_22(MultLoop_acc_694_itm_19_2_1) +
      ({(data_rsci_idat[71:54]) , 4'b0001});
  assign MultLoop_acc_1380_nl = nl_MultLoop_acc_1380_nl[21:0];
  assign nl_MultLoop_acc_972_nl = ({(data_rsci_idat[107:90]) , 2'b01}) + conv_s2s_19_20({Result_Result_conc_60_18_7
      , (~ (data_rsci_idat[96:90]))});
  assign MultLoop_acc_972_nl = nl_MultLoop_acc_972_nl[19:0];
  assign nl_MultLoop_acc_973_nl = ({(~ (data_rsci_idat[107:90])) , 4'b0000}) + conv_s2s_20_22(MultLoop_acc_972_nl);
  assign MultLoop_acc_973_nl = nl_MultLoop_acc_973_nl[21:0];
  assign nl_MultLoop_acc_82_nl = conv_s2s_22_26(MultLoop_acc_973_nl) + conv_s2s_25_26({(~
      (data_rsci_idat[107:90])) , 7'b0010000});
  assign MultLoop_acc_82_nl = nl_MultLoop_acc_82_nl[25:0];
  assign nl_MultLoop_acc_966_nl = ({(~ (data_rsci_idat[17:0])) , 4'b0000}) + conv_s2s_20_22(MultLoop_acc_805_cse_1);
  assign MultLoop_acc_966_nl = nl_MultLoop_acc_966_nl[21:0];
  assign nl_MultLoop_acc_77_nl = conv_s2s_22_24(MultLoop_acc_966_nl) + ({(data_rsci_idat[17:0])
      , 6'b010000});
  assign MultLoop_acc_77_nl = nl_MultLoop_acc_77_nl[23:0];
  assign nl_MultLoop_acc_1297_nl =  -conv_s2s_14_15(data_rsci_idat[35:22]);
  assign MultLoop_acc_1297_nl = nl_MultLoop_acc_1297_nl[14:0];
  assign nl_MultLoop_acc_964_nl = ({(data_rsci_idat[35:18]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_1297_nl)
      , (~ (data_rsci_idat[21:18]))});
  assign MultLoop_acc_964_nl = nl_MultLoop_acc_964_nl[19:0];
  assign nl_MultLoop_acc_78_nl = conv_s2s_20_22(MultLoop_acc_964_nl) + ({(~ (data_rsci_idat[35:18]))
      , 4'b0000});
  assign MultLoop_acc_78_nl = nl_MultLoop_acc_78_nl[21:0];
  assign nl_MultLoop_acc_984_nl = (readslicef_26_16_10((MultLoop_acc_82_nl))) + conv_s2s_14_16(readslicef_24_14_10((MultLoop_acc_77_nl)))
      + conv_s2s_12_16(readslicef_22_12_10((MultLoop_acc_78_nl))) + 16'b1111111001111001;
  assign MultLoop_acc_984_nl = nl_MultLoop_acc_984_nl[15:0];
  assign nl_MultLoop_acc_986_nl = conv_s2s_17_18(readslicef_22_17_5((MultLoop_acc_1380_nl)))
      + conv_s2s_16_18(MultLoop_acc_984_nl);
  assign MultLoop_acc_986_nl = nl_MultLoop_acc_986_nl[17:0];
  assign nl_MultLoop_acc_989_nl = (MultLoop_acc_986_nl) + MultLoop_acc_1374_itm_18_1;
  assign MultLoop_acc_989_nl = nl_MultLoop_acc_989_nl[17:0];
  assign nl_MultLoop_acc_975_nl = conv_s2s_18_19(data_rsci_idat[179:162]) + conv_s2s_17_19({MultLoop_MultLoop_conc_226_16_4
      , (data_rsci_idat[167:164])});
  assign MultLoop_acc_975_nl = nl_MultLoop_acc_975_nl[18:0];
  assign nl_MultLoop_acc_86_nl = conv_s2u_19_22(MultLoop_acc_975_nl) + ({(~ (data_rsci_idat[179:162]))
      , 4'b0000});
  assign MultLoop_acc_86_nl = nl_MultLoop_acc_86_nl[21:0];
  assign nl_MultLoop_acc_1293_nl = conv_s2u_13_18(MultLoop_acc_916_itm_18_3[15:3])
      + (~ (data_rsci_idat[143:126]));
  assign MultLoop_acc_1293_nl = nl_MultLoop_acc_1293_nl[17:0];
  assign nl_MultLoop_acc_969_nl = (~ (data_rsci_idat[89:72])) + conv_s2s_14_18(data_rsci_idat[89:76]);
  assign MultLoop_acc_969_nl = nl_MultLoop_acc_969_nl[17:0];
  assign nl_MultLoop_acc_970_nl = conv_s2s_20_21({(~ (data_rsci_idat[89:72])) , 2'b01})
      + conv_s2s_18_21(MultLoop_acc_969_nl);
  assign MultLoop_acc_970_nl = nl_MultLoop_acc_970_nl[20:0];
  assign nl_MultLoop_acc_315_nl = conv_s2u_21_22(MultLoop_acc_970_nl) + ({(data_rsci_idat[89:72])
      , 4'b0100});
  assign MultLoop_acc_315_nl = nl_MultLoop_acc_315_nl[21:0];
  assign nl_MultLoop_acc_976_nl = conv_s2s_21_22({(~ (data_rsci_idat[125:108])) ,
      3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[125:108]));
  assign MultLoop_acc_976_nl = nl_MultLoop_acc_976_nl[21:0];
  assign nl_MultLoop_acc_83_nl = conv_s2s_22_27(MultLoop_acc_976_nl) + ({(data_rsci_idat[125:108])
      , 9'b000001000});
  assign MultLoop_acc_83_nl = nl_MultLoop_acc_83_nl[26:0];
  assign nl_MultLoop_acc_1295_nl =  -conv_s2s_14_15(data_rsci_idat[53:40]);
  assign MultLoop_acc_1295_nl = nl_MultLoop_acc_1295_nl[14:0];
  assign nl_MultLoop_acc_79_nl = conv_s2s_22_23({(~ (data_rsci_idat[53:36])) , 4'b0100})
      + conv_s2s_20_23({(~ (data_rsci_idat[53:36])) , 2'b01}) + conv_s2s_19_23({(MultLoop_acc_1295_nl)
      , (~ (data_rsci_idat[39:36]))});
  assign MultLoop_acc_79_nl = nl_MultLoop_acc_79_nl[22:0];
  assign nl_res_rsci_d_125_108  = (MultLoop_acc_989_nl) + conv_s2s_17_18(readslicef_22_17_5((MultLoop_acc_86_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_1293_nl))) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_315_nl)))
      + conv_s2s_17_18(readslicef_27_17_10((MultLoop_acc_83_nl))) + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_79_nl)));
  assign nl_MultLoop_acc_496_nl = ({(data_rsci_idat[143:126]) , 6'b010000}) + conv_s2s_22_24({(~
      (data_rsci_idat[143:126])) , 4'b0100}) + conv_s2s_21_24(MultLoop_acc_406_cse_1);
  assign MultLoop_acc_496_nl = nl_MultLoop_acc_496_nl[23:0];
  assign nl_MultLoop_acc_1287_nl = conv_s2u_16_19(readslicef_24_16_8((MultLoop_acc_496_nl)))
      + conv_s2u_18_19(data_rsci_idat[143:126]);
  assign MultLoop_acc_1287_nl = nl_MultLoop_acc_1287_nl[18:0];
  assign nl_MultLoop_acc_501_nl = conv_s2s_13_14(MultLoop_acc_237_itm_22_9[13:1])
      + 14'b00001101110011;
  assign MultLoop_acc_501_nl = nl_MultLoop_acc_501_nl[13:0];
  assign nl_MultLoop_acc_499_nl = ({(data_rsci_idat[35:18]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[35:18])) , 2'b01}) + conv_s2s_19_22({MultLoop_MultLoop_conc_210_18_8
      , (~ (data_rsci_idat[25:18]))});
  assign MultLoop_acc_499_nl = nl_MultLoop_acc_499_nl[21:0];
  assign nl_MultLoop_acc_1289_nl = (~ (data_rsci_idat[35:18])) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_499_nl)));
  assign MultLoop_acc_1289_nl = nl_MultLoop_acc_1289_nl[17:0];
  assign nl_MultLoop_acc_1290_nl = conv_s2u_18_21(MultLoop_acc_1289_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[35:18])) , 2'b01});
  assign MultLoop_acc_1290_nl = nl_MultLoop_acc_1290_nl[20:0];
  assign nl_MultLoop_242_MultLoop_acc_3_nl = conv_s2s_14_17(MultLoop_acc_501_nl)
      + (readslicef_21_17_4((MultLoop_acc_1290_nl)));
  assign MultLoop_242_MultLoop_acc_3_nl = nl_MultLoop_242_MultLoop_acc_3_nl[16:0];
  assign nl_MultLoop_acc_1291_nl =  -conv_s2s_16_17(data_rsci_idat[71:56]);
  assign MultLoop_acc_1291_nl = nl_MultLoop_acc_1291_nl[16:0];
  assign nl_MultLoop_acc_270_nl = conv_s2s_19_21({(MultLoop_acc_1291_nl) , (~ (data_rsci_idat[55:54]))})
      + conv_s2s_20_21({(~ (data_rsci_idat[71:54])) , 2'b01});
  assign MultLoop_acc_270_nl = nl_MultLoop_acc_270_nl[20:0];
  assign nl_MultLoop_acc_1379_nl = conv_s2u_19_24(MultLoop_acc_808_itm_20_2_1) +
      ({(data_rsci_idat[125:108]) , 6'b000001});
  assign MultLoop_acc_1379_nl = nl_MultLoop_acc_1379_nl[23:0];
  assign nl_MultLoop_acc_510_nl = conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_1287_nl)))
      + conv_s2s_17_18(MultLoop_242_MultLoop_acc_3_nl) + conv_s2s_17_18(readslicef_21_17_4((MultLoop_acc_270_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1379_nl)));
  assign MultLoop_acc_510_nl = nl_MultLoop_acc_510_nl[17:0];
  assign nl_MultLoop_acc_1282_nl = conv_s2s_14_15(data_rsci_idat[53:40]) + 15'b000000000000001;
  assign MultLoop_acc_1282_nl = nl_MultLoop_acc_1282_nl[14:0];
  assign nl_MultLoop_acc_504_nl = conv_s2s_18_19(data_rsci_idat[53:36]) + conv_s2s_17_19({(MultLoop_acc_1282_nl)
      , (data_rsci_idat[39:38])});
  assign MultLoop_acc_504_nl = nl_MultLoop_acc_504_nl[18:0];
  assign nl_MultLoop_acc_269_nl = conv_s2u_19_20(MultLoop_acc_504_nl) + ({(~ (data_rsci_idat[53:36]))
      , 2'b00});
  assign MultLoop_acc_269_nl = nl_MultLoop_acc_269_nl[19:0];
  assign nl_MultLoop_acc_1393_nl = conv_s2u_18_19(data_rsci_idat[107:90]) + conv_s2u_17_19(MultLoop_acc_753_cse_1[18:2]);
  assign MultLoop_acc_1393_nl = nl_MultLoop_acc_1393_nl[18:0];
  assign nl_MultLoop_acc_1284_nl = conv_s2u_15_18(readslicef_19_15_4((MultLoop_acc_1393_nl)))
      + (~ (data_rsci_idat[107:90]));
  assign MultLoop_acc_1284_nl = nl_MultLoop_acc_1284_nl[17:0];
  assign nl_MultLoop_acc_485_nl = ({(~ (data_rsci_idat[89:72])) , 4'b0000}) + conv_s2s_20_22(MultLoop_acc_786_cse_1);
  assign MultLoop_acc_485_nl = nl_MultLoop_acc_485_nl[21:0];
  assign nl_MultLoop_acc_271_nl = conv_s2s_22_25(MultLoop_acc_485_nl) + ({(data_rsci_idat[89:72])
      , 7'b0010000});
  assign MultLoop_acc_271_nl = nl_MultLoop_acc_271_nl[24:0];
  assign nl_MultLoop_acc_505_nl = conv_s2s_16_17(readslicef_18_16_2((MultLoop_acc_1284_nl)))
      + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_271_nl)));
  assign MultLoop_acc_505_nl = nl_MultLoop_acc_505_nl[16:0];
  assign nl_MultLoop_acc_509_nl = (readslicef_20_18_2((MultLoop_acc_269_nl))) + conv_s2s_17_18(MultLoop_acc_505_nl);
  assign MultLoop_acc_509_nl = nl_MultLoop_acc_509_nl[17:0];
  assign nl_MultLoop_acc_490_nl = conv_s2s_18_19(data_rsci_idat[161:144]) + conv_s2s_14_19(data_rsci_idat[161:148]);
  assign MultLoop_acc_490_nl = nl_MultLoop_acc_490_nl[18:0];
  assign nl_MultLoop_acc_365_nl = conv_s2u_19_21(MultLoop_acc_490_nl) + conv_s2u_20_21({(data_rsci_idat[161:144])
      , 2'b00});
  assign MultLoop_acc_365_nl = nl_MultLoop_acc_365_nl[20:0];
  assign nl_MultLoop_acc_492_nl = (~ (data_rsci_idat[179:162])) + conv_s2s_17_18({MultLoop_MultLoop_conc_224_16_6
      , (data_rsci_idat[169:164])});
  assign MultLoop_acc_492_nl = nl_MultLoop_acc_492_nl[17:0];
  assign nl_MultLoop_acc_493_nl = ({(data_rsci_idat[179:162]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_492_nl);
  assign MultLoop_acc_493_nl = nl_MultLoop_acc_493_nl[19:0];
  assign nl_MultLoop_acc_1286_nl = conv_s2u_14_18(readslicef_20_14_6((MultLoop_acc_493_nl)))
      + (~ (data_rsci_idat[179:162]));
  assign MultLoop_acc_1286_nl = nl_MultLoop_acc_1286_nl[17:0];
  assign nl_res_rsci_d_449_432  = (MultLoop_acc_510_nl) + (MultLoop_acc_509_nl) +
      conv_s2s_17_18(readslicef_21_17_4((MultLoop_acc_365_nl))) + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_1286_nl)));
  assign nl_MultLoop_acc_1278_nl =  -conv_s2s_10_11(data_rsci_idat[143:134]);
  assign MultLoop_acc_1278_nl = nl_MultLoop_acc_1278_nl[10:0];
  assign nl_MultLoop_acc_95_nl = conv_s2s_19_27({(MultLoop_acc_1278_nl) , (~ (data_rsci_idat[133:126]))})
      + conv_s2s_26_27({(~ (data_rsci_idat[143:126])) , 8'b00000001});
  assign MultLoop_acc_95_nl = nl_MultLoop_acc_95_nl[26:0];
  assign nl_MultLoop_acc_1279_nl =  -conv_s2s_9_10(data_rsci_idat[53:45]);
  assign MultLoop_acc_1279_nl = nl_MultLoop_acc_1279_nl[9:0];
  assign nl_MultLoop_acc_947_nl = ({(data_rsci_idat[53:36]) , 5'b01000}) + conv_s2s_21_23({(~
      (data_rsci_idat[53:36])) , 3'b001}) + conv_s2s_19_23({(MultLoop_acc_1279_nl)
      , (~ (data_rsci_idat[44:36]))});
  assign MultLoop_acc_947_nl = nl_MultLoop_acc_947_nl[22:0];
  assign nl_MultLoop_acc_1280_nl = conv_s2u_18_19(data_rsci_idat[53:36]) + conv_s2u_16_19(readslicef_23_16_7((MultLoop_acc_947_nl)));
  assign MultLoop_acc_1280_nl = nl_MultLoop_acc_1280_nl[18:0];
  assign nl_MultLoop_acc_1281_nl = conv_s2u_17_18(readslicef_19_17_2((MultLoop_acc_1280_nl)))
      + (~ (data_rsci_idat[53:36]));
  assign MultLoop_acc_1281_nl = nl_MultLoop_acc_1281_nl[17:0];
  assign nl_MultLoop_71_MultLoop_acc_3_nl = nnet_product_input_t_config2_weight_t_config2_accum_t_acc_4_itm_18_2_1
      + 17'b00000000111100101;
  assign MultLoop_71_MultLoop_acc_3_nl = nl_MultLoop_71_MultLoop_acc_3_nl[16:0];
  assign nl_MultLoop_acc_961_nl = conv_s2s_17_18(readslicef_27_17_10((MultLoop_acc_95_nl)))
      + conv_s2s_17_18(MultLoop_acc_1354_itm_19_3) + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_1281_nl)))
      + conv_s2s_17_18(MultLoop_71_MultLoop_acc_3_nl);
  assign MultLoop_acc_961_nl = nl_MultLoop_acc_961_nl[17:0];
  assign nl_MultLoop_acc_1377_nl = conv_s2u_15_19(MultLoop_acc_812_cse_1[18:4]) +
      conv_s2u_18_19(data_rsci_idat[35:18]);
  assign MultLoop_acc_1377_nl = nl_MultLoop_acc_1377_nl[18:0];
  assign nl_MultLoop_acc_317_nl = conv_s2u_18_21(MultLoop_acc_621_cse_1) + ({(data_rsci_idat[125:108])
      , 3'b001});
  assign MultLoop_acc_317_nl = nl_MultLoop_acc_317_nl[20:0];
  assign nl_MultLoop_acc_956_nl = conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_1377_nl)))
      + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_317_nl)));
  assign MultLoop_acc_956_nl = nl_MultLoop_acc_956_nl[17:0];
  assign nl_MultLoop_acc_950_nl = (~ (data_rsci_idat[161:144])) + conv_s2s_15_18(data_rsci_idat[161:147]);
  assign MultLoop_acc_950_nl = nl_MultLoop_acc_950_nl[17:0];
  assign nl_MultLoop_acc_951_nl = ({(data_rsci_idat[161:144]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_950_nl);
  assign MultLoop_acc_951_nl = nl_MultLoop_acc_951_nl[19:0];
  assign nl_MultLoop_acc_318_nl = conv_s2u_20_24(MultLoop_acc_951_nl) + conv_s2u_23_24({(data_rsci_idat[161:144])
      , 5'b00000});
  assign MultLoop_acc_318_nl = nl_MultLoop_acc_318_nl[23:0];
  assign nl_MultLoop_acc_960_nl = (MultLoop_acc_956_nl) + (readslicef_24_18_6((MultLoop_acc_318_nl)));
  assign MultLoop_acc_960_nl = nl_MultLoop_acc_960_nl[17:0];
  assign nl_MultLoop_acc_954_nl = conv_s2s_20_21({(data_rsci_idat[179:162]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[179:162]) + conv_s2s_17_21({MultLoop_acc_1273_cse_1
      , (data_rsci_idat[170:164])});
  assign MultLoop_acc_954_nl = nl_MultLoop_acc_954_nl[20:0];
  assign nl_MultLoop_acc_1274_nl = conv_s2u_14_18(readslicef_21_14_7((MultLoop_acc_954_nl)))
      + (~ (data_rsci_idat[179:162]));
  assign MultLoop_acc_1274_nl = nl_MultLoop_acc_1274_nl[17:0];
  assign nl_MultLoop_acc_1275_nl = conv_s2s_12_13(data_rsci_idat[107:96]) + 13'b0000000000001;
  assign MultLoop_acc_1275_nl = nl_MultLoop_acc_1275_nl[12:0];
  assign nl_MultLoop_acc_942_nl = conv_s2s_18_19(data_rsci_idat[107:90]) + conv_s2s_15_19({(MultLoop_acc_1275_nl)
      , (data_rsci_idat[95:94])});
  assign MultLoop_acc_942_nl = nl_MultLoop_acc_942_nl[18:0];
  assign nl_MultLoop_acc_93_nl = conv_s2u_19_20(MultLoop_acc_942_nl) + ({(~ (data_rsci_idat[107:90]))
      , 2'b00});
  assign MultLoop_acc_93_nl = nl_MultLoop_acc_93_nl[19:0];
  assign nl_MultLoop_acc_1411_nl = ({(data_rsci_idat[71:54]) , 2'b01}) + conv_s2u_19_20(MultLoop_acc_1397_itm_21_3_1);
  assign MultLoop_acc_1411_nl = nl_MultLoop_acc_1411_nl[19:0];
  assign nl_MultLoop_acc_1277_nl = conv_s2u_16_18(readslicef_20_16_4((MultLoop_acc_1411_nl)))
      + (~ (data_rsci_idat[71:54]));
  assign MultLoop_acc_1277_nl = nl_MultLoop_acc_1277_nl[17:0];
  assign nl_MultLoop_acc_955_nl = conv_s2s_16_17(readslicef_20_16_4((MultLoop_acc_93_nl)))
      + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_1277_nl)));
  assign MultLoop_acc_955_nl = nl_MultLoop_acc_955_nl[16:0];
  assign nl_MultLoop_acc_959_nl = (MultLoop_acc_1274_nl) + conv_s2s_17_18(MultLoop_acc_955_nl);
  assign MultLoop_acc_959_nl = nl_MultLoop_acc_959_nl[17:0];
  assign nl_res_rsci_d_143_126  = (MultLoop_acc_961_nl) + (MultLoop_acc_960_nl) +
      (MultLoop_acc_959_nl);
  assign nl_MultLoop_acc_525_nl = conv_s2s_23_24({(~ (data_rsci_idat[53:36])) , 5'b01000})
      + conv_s2s_22_24(MultLoop_acc_560_cse_1);
  assign MultLoop_acc_525_nl = nl_MultLoop_acc_525_nl[23:0];
  assign nl_MultLoop_acc_260_nl = conv_s2s_24_25(MultLoop_acc_525_nl) + ({(data_rsci_idat[53:36])
      , 7'b0100000});
  assign MultLoop_acc_260_nl = nl_MultLoop_acc_260_nl[24:0];
  assign nl_MultLoop_acc_521_nl = conv_s2s_23_24({(~ (data_rsci_idat[107:90])) ,
      5'b01000}) + conv_s2s_21_24({(~ (data_rsci_idat[107:90])) , 3'b001}) + conv_s2s_18_24(~
      (data_rsci_idat[107:90]));
  assign MultLoop_acc_521_nl = nl_MultLoop_acc_521_nl[23:0];
  assign nl_MultLoop_acc_263_nl = conv_s2s_24_26(MultLoop_acc_521_nl) + ({(data_rsci_idat[107:90])
      , 8'b00100000});
  assign MultLoop_acc_263_nl = nl_MultLoop_acc_263_nl[25:0];
  assign nl_MultLoop_acc_1406_nl = conv_s2u_19_23(MultLoop_acc_1397_itm_21_3_1) +
      conv_s2u_22_23({(~ (data_rsci_idat[71:54])) , 4'b0001});
  assign MultLoop_acc_1406_nl = nl_MultLoop_acc_1406_nl[22:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_13_nl = (readslicef_25_18_7((MultLoop_acc_260_nl)))
      + conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_263_nl))) + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_1406_nl)));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_13_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_13_nl[17:0];
  assign nl_MultLoop_acc_526_nl = ({(data_rsci_idat[179:162]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[179:162]));
  assign MultLoop_acc_526_nl = nl_MultLoop_acc_526_nl[20:0];
  assign nl_MultLoop_acc_1267_nl = (~ (data_rsci_idat[179:162])) + conv_s2s_15_18(readslicef_21_15_6((MultLoop_acc_526_nl)));
  assign MultLoop_acc_1267_nl = nl_MultLoop_acc_1267_nl[17:0];
  assign nl_MultLoop_acc_1268_nl = conv_s2u_18_21(MultLoop_acc_1267_nl) + ({(data_rsci_idat[179:162])
      , 3'b001});
  assign MultLoop_acc_1268_nl = nl_MultLoop_acc_1268_nl[20:0];
  assign nl_MultLoop_acc_1269_nl = conv_s2s_12_13(data_rsci_idat[35:24]) + 13'b0000000000001;
  assign MultLoop_acc_1269_nl = nl_MultLoop_acc_1269_nl[12:0];
  assign nl_MultLoop_acc_513_nl = conv_s2s_18_19(data_rsci_idat[35:18]) + conv_s2s_17_19({(MultLoop_acc_1269_nl)
      , (data_rsci_idat[23:20])});
  assign MultLoop_acc_513_nl = nl_MultLoop_acc_513_nl[18:0];
  assign nl_MultLoop_acc_259_nl = conv_s2u_19_22(MultLoop_acc_513_nl) + ({(~ (data_rsci_idat[35:18]))
      , 4'b0000});
  assign MultLoop_acc_259_nl = nl_MultLoop_acc_259_nl[21:0];
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_nor_nl = ~((data_rsci_idat[146:144]!=3'b000));
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_7_nl = conv_s2s_15_16(~
      (data_rsci_idat[161:147])) + conv_s2s_14_16(readslicef_22_14_8((MultLoop_acc_259_nl)))
      + conv_u2s_1_16(nnet_product_input_t_config2_weight_t_config2_accum_t_nor_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_7_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_7_nl[15:0];
  assign nl_MultLoop_acc_515_nl = conv_s2s_21_22({(data_rsci_idat[125:108]) , 3'b000})
      + conv_s2s_19_22(MultLoop_acc_650_cse_1);
  assign MultLoop_acc_515_nl = nl_MultLoop_acc_515_nl[21:0];
  assign nl_MultLoop_acc_364_nl = conv_s2u_22_24(MultLoop_acc_515_nl) + conv_s2u_23_24({(data_rsci_idat[125:108])
      , 5'b00000});
  assign MultLoop_acc_364_nl = nl_MultLoop_acc_364_nl[23:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_9_nl = conv_s2s_16_17(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_7_nl)
      + conv_s2s_16_17(readslicef_24_16_8((MultLoop_acc_364_nl)));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_9_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_9_nl[16:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_12_nl = (readslicef_21_18_3((MultLoop_acc_1268_nl)))
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_9_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_12_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_12_nl[17:0];
  assign nl_MultLoop_acc_1270_nl =  -conv_s2s_12_13(data_rsci_idat[143:132]);
  assign MultLoop_acc_1270_nl = nl_MultLoop_acc_1270_nl[12:0];
  assign nl_MultLoop_acc_519_nl = ({(data_rsci_idat[143:126]) , 4'b0001}) + conv_s2s_19_22({(MultLoop_acc_1270_nl)
      , (~ (data_rsci_idat[131:126]))});
  assign MultLoop_acc_519_nl = nl_MultLoop_acc_519_nl[21:0];
  assign nl_MultLoop_acc_1271_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_519_nl)))
      + (~ (data_rsci_idat[143:126]));
  assign MultLoop_acc_1271_nl = nl_MultLoop_acc_1271_nl[17:0];
  assign nl_MultLoop_acc_1376_nl = conv_s2u_19_21(MultLoop_acc_399_cse_1[20:2]) +
      ({(data_rsci_idat[17:0]) , 3'b001});
  assign MultLoop_acc_1376_nl = nl_MultLoop_acc_1376_nl[20:0];
  assign nl_MultLoop_231_MultLoop_acc_3_nl = (readslicef_21_16_5((MultLoop_acc_1376_nl)))
      + 16'b1111111011100001;
  assign MultLoop_231_MultLoop_acc_3_nl = nl_MultLoop_231_MultLoop_acc_3_nl[15:0];
  assign nl_res_rsci_d_431_414  = (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_13_nl)
      + (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_12_nl) + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_1271_nl)))
      + conv_s2s_16_18(MultLoop_acc_114_itm_19_3[16:1]) + conv_s2s_16_18(MultLoop_231_MultLoop_acc_3_nl);
  assign nl_MultLoop_acc_925_nl = conv_s2s_24_25({(~ (data_rsci_idat[89:72])) , 6'b010000})
      + conv_s2s_22_25({(~ (data_rsci_idat[89:72])) , 4'b0100}) + conv_s2s_21_25(MultLoop_acc_745_cse_1);
  assign MultLoop_acc_925_nl = nl_MultLoop_acc_925_nl[24:0];
  assign nl_MultLoop_acc_104_nl = conv_s2s_25_26(MultLoop_acc_925_nl) + ({(data_rsci_idat[89:72])
      , 8'b01000000});
  assign MultLoop_acc_104_nl = nl_MultLoop_acc_104_nl[25:0];
  assign nl_MultLoop_acc_99_nl = (MultLoop_acc_100_itm_23_7[16:2]) + 15'b000000000000001;
  assign MultLoop_acc_99_nl = nl_MultLoop_acc_99_nl[14:0];
  assign nl_MultLoop_acc_1392_nl = conv_s2u_18_19(data_rsci_idat[143:126]) + conv_s2u_16_19(MultLoop_acc_916_itm_18_3);
  assign MultLoop_acc_1392_nl = nl_MultLoop_acc_1392_nl[18:0];
  assign nl_MultLoop_acc_1266_nl = conv_s2u_16_18(readslicef_19_16_3((MultLoop_acc_1392_nl)))
      + (~ (data_rsci_idat[143:126]));
  assign MultLoop_acc_1266_nl = nl_MultLoop_acc_1266_nl[17:0];
  assign nl_MultLoop_acc_935_nl = (readslicef_26_18_8((MultLoop_acc_104_nl))) + conv_s2s_17_18({(MultLoop_acc_99_nl)
      , (MultLoop_acc_100_itm_23_7[1:0])}) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_1266_nl)));
  assign MultLoop_acc_935_nl = nl_MultLoop_acc_935_nl[17:0];
  assign nl_MultLoop_acc_927_nl = ({(~ (data_rsci_idat[179:162])) , 4'b0000}) + conv_s2s_19_22(MultLoop_acc_702_cse_1);
  assign MultLoop_acc_927_nl = nl_MultLoop_acc_927_nl[21:0];
  assign nl_MultLoop_acc_928_nl = conv_s2s_24_25({(~ (data_rsci_idat[179:162])) ,
      6'b010000}) + conv_s2s_22_25(MultLoop_acc_927_nl);
  assign MultLoop_acc_928_nl = nl_MultLoop_acc_928_nl[24:0];
  assign nl_MultLoop_acc_321_nl = conv_s2u_25_26(MultLoop_acc_928_nl) + ({(data_rsci_idat[179:162])
      , 8'b01000000});
  assign MultLoop_acc_321_nl = nl_MultLoop_acc_321_nl[25:0];
  assign nl_MultLoop_acc_918_nl = conv_s2s_18_19(data_rsci_idat[107:90]) + conv_s2s_15_19(data_rsci_idat[107:93]);
  assign MultLoop_acc_918_nl = nl_MultLoop_acc_918_nl[18:0];
  assign nl_MultLoop_acc_320_nl = conv_s2u_19_23(MultLoop_acc_918_nl) + conv_s2u_22_23({(data_rsci_idat[107:90])
      , 4'b0000});
  assign MultLoop_acc_320_nl = nl_MultLoop_acc_320_nl[22:0];
  assign nl_MultLoop_acc_919_nl = ({(data_rsci_idat[71:54]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[71:54]));
  assign MultLoop_acc_919_nl = nl_MultLoop_acc_919_nl[19:0];
  assign nl_MultLoop_acc_103_nl = conv_s2s_24_25({(data_rsci_idat[71:54]) , 6'b000000})
      + conv_s2s_22_25({(data_rsci_idat[71:54]) , 4'b0000}) + conv_s2s_20_25(MultLoop_acc_919_nl);
  assign MultLoop_acc_103_nl = nl_MultLoop_acc_103_nl[24:0];
  assign nl_MultLoop_acc_931_nl = conv_s2s_16_17(readslicef_23_16_7((MultLoop_acc_320_nl)))
      + conv_s2s_16_17(readslicef_25_16_9((MultLoop_acc_103_nl)));
  assign MultLoop_acc_931_nl = nl_MultLoop_acc_931_nl[16:0];
  assign nl_MultLoop_acc_934_nl = (readslicef_26_18_8((MultLoop_acc_321_nl))) + conv_s2s_17_18(MultLoop_acc_931_nl);
  assign MultLoop_acc_934_nl = nl_MultLoop_acc_934_nl[17:0];
  assign nl_MultLoop_acc_922_nl = ({(data_rsci_idat[125:108]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[125:108]));
  assign MultLoop_acc_922_nl = nl_MultLoop_acc_922_nl[19:0];
  assign nl_MultLoop_acc_1264_nl = conv_s2u_12_19(readslicef_20_12_8((MultLoop_acc_922_nl)))
      + conv_s2u_18_19(data_rsci_idat[125:108]);
  assign MultLoop_acc_1264_nl = nl_MultLoop_acc_1264_nl[18:0];
  assign nl_MultLoop_acc_921_nl = conv_s2s_22_23({(~ (data_rsci_idat[35:18])) , 4'b0001})
      + conv_s2s_18_23(~ (data_rsci_idat[35:18]));
  assign MultLoop_acc_921_nl = nl_MultLoop_acc_921_nl[22:0];
  assign nl_MultLoop_acc_101_nl = conv_s2s_23_25(MultLoop_acc_921_nl) + ({(data_rsci_idat[35:18])
      , 7'b0010000});
  assign MultLoop_acc_101_nl = nl_MultLoop_acc_101_nl[24:0];
  assign nl_MultLoop_acc_914_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_15_18(data_rsci_idat[53:39]);
  assign MultLoop_acc_914_nl = nl_MultLoop_acc_914_nl[17:0];
  assign nl_MultLoop_acc_319_nl = conv_s2u_18_20(MultLoop_acc_914_nl) + ({(data_rsci_idat[53:36])
      , 2'b01});
  assign MultLoop_acc_319_nl = nl_MultLoop_acc_319_nl[19:0];
  assign nl_res_rsci_d_161_144  = (MultLoop_acc_935_nl) + (MultLoop_acc_934_nl) +
      conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_1264_nl))) + conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_101_nl)))
      + conv_s2s_13_18(MultLoop_acc_108_itm_19_6[13:1]) + conv_s2s_13_18(readslicef_20_13_7((MultLoop_acc_319_nl)));
  assign nl_MultLoop_acc_542_nl = (~ (data_rsci_idat[17:0])) + conv_s2s_16_18({MultLoop_acc_1239_cse_1
      , (data_rsci_idat[4:3])});
  assign MultLoop_acc_542_nl = nl_MultLoop_acc_542_nl[17:0];
  assign nl_MultLoop_acc_360_nl = conv_s2u_18_21(MultLoop_acc_542_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[17:0])) , 2'b01});
  assign MultLoop_acc_360_nl = nl_MultLoop_acc_360_nl[20:0];
  assign nl_MultLoop_acc_544_nl = ({(data_rsci_idat[35:18]) , 4'b0001}) + conv_s2s_18_22(MultLoop_acc_543_cse_1);
  assign MultLoop_acc_544_nl = nl_MultLoop_acc_544_nl[21:0];
  assign nl_MultLoop_acc_1256_nl = conv_s2u_15_19(readslicef_22_15_7((MultLoop_acc_544_nl)))
      + conv_s2u_18_19(data_rsci_idat[35:18]);
  assign MultLoop_acc_1256_nl = nl_MultLoop_acc_1256_nl[18:0];
  assign nl_MultLoop_acc_551_nl = (readslicef_21_18_3((MultLoop_acc_360_nl))) + (readslicef_19_18_1((MultLoop_acc_1256_nl)));
  assign MultLoop_acc_551_nl = nl_MultLoop_acc_551_nl[17:0];
  assign nl_MultLoop_acc_529_nl = conv_s2s_21_22({(~ (data_rsci_idat[143:126])) ,
      3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[143:126]));
  assign MultLoop_acc_529_nl = nl_MultLoop_acc_529_nl[21:0];
  assign nl_MultLoop_acc_254_nl = conv_s2s_22_23(MultLoop_acc_529_nl) + ({(data_rsci_idat[143:126])
      , 5'b01000});
  assign MultLoop_acc_254_nl = nl_MultLoop_acc_254_nl[22:0];
  assign nl_MultLoop_acc_531_nl = ({(data_rsci_idat[53:36]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_218_18_8
      , (~ (data_rsci_idat[43:36]))});
  assign MultLoop_acc_531_nl = nl_MultLoop_acc_531_nl[19:0];
  assign nl_MultLoop_acc_532_nl = conv_s2s_22_23({(data_rsci_idat[53:36]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_531_nl);
  assign MultLoop_acc_532_nl = nl_MultLoop_acc_532_nl[22:0];
  assign nl_MultLoop_acc_1258_nl = conv_s2u_15_18(readslicef_23_15_8((MultLoop_acc_532_nl)))
      + (~ (data_rsci_idat[53:36]));
  assign MultLoop_acc_1258_nl = nl_MultLoop_acc_1258_nl[17:0];
  assign nl_MultLoop_acc_362_nl = conv_s2u_15_19(data_rsci_idat[71:57]) + conv_s2u_18_19(data_rsci_idat[71:54]);
  assign MultLoop_acc_362_nl = nl_MultLoop_acc_362_nl[18:0];
  assign nl_MultLoop_acc_1259_nl =  -conv_s2s_15_16(data_rsci_idat[125:111]);
  assign MultLoop_acc_1259_nl = nl_MultLoop_acc_1259_nl[15:0];
  assign nl_MultLoop_acc_253_nl = conv_s2s_19_22({(MultLoop_acc_1259_nl) , (~ (data_rsci_idat[110:108]))})
      + conv_s2s_21_22({(~ (data_rsci_idat[125:108])) , 3'b001});
  assign MultLoop_acc_253_nl = nl_MultLoop_acc_253_nl[21:0];
  assign nl_MultLoop_acc_545_nl = (readslicef_22_13_9((MultLoop_acc_253_nl))) + 13'b0000000110111;
  assign MultLoop_acc_545_nl = nl_MultLoop_acc_545_nl[12:0];
  assign nl_MultLoop_acc_550_nl = conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_254_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_1258_nl))) + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_362_nl)))
      + conv_s2s_13_18(MultLoop_acc_545_nl);
  assign MultLoop_acc_550_nl = nl_MultLoop_acc_550_nl[17:0];
  assign nl_MultLoop_acc_553_nl = (MultLoop_acc_551_nl) + (MultLoop_acc_550_nl);
  assign MultLoop_acc_553_nl = nl_MultLoop_acc_553_nl[17:0];
  assign nl_MultLoop_acc_533_nl = (~ (data_rsci_idat[179:162])) + conv_s2s_15_18(data_rsci_idat[179:165]);
  assign MultLoop_acc_533_nl = nl_MultLoop_acc_533_nl[17:0];
  assign nl_MultLoop_acc_534_nl = conv_s2s_20_21({(~ (data_rsci_idat[179:162])) ,
      2'b01}) + conv_s2s_18_21(MultLoop_acc_533_nl);
  assign MultLoop_acc_534_nl = nl_MultLoop_acc_534_nl[20:0];
  assign nl_MultLoop_acc_363_nl = conv_s2u_21_22(MultLoop_acc_534_nl) + ({(data_rsci_idat[179:162])
      , 4'b0100});
  assign MultLoop_acc_363_nl = nl_MultLoop_acc_363_nl[21:0];
  assign nl_MultLoop_acc_1410_nl = conv_s2u_18_19(data_rsci_idat[89:72]) + conv_s2u_16_19(MultLoop_acc_1399_itm_20_5);
  assign MultLoop_acc_1410_nl = nl_MultLoop_acc_1410_nl[18:0];
  assign nl_MultLoop_acc_1261_nl = conv_s2u_18_19(data_rsci_idat[89:72]) + conv_s2u_17_19(readslicef_19_17_2((MultLoop_acc_1410_nl)));
  assign MultLoop_acc_1261_nl = nl_MultLoop_acc_1261_nl[18:0];
  assign nl_MultLoop_acc_1262_nl = conv_s2u_17_18(readslicef_19_17_2((MultLoop_acc_1261_nl)))
      + (~ (data_rsci_idat[89:72]));
  assign MultLoop_acc_1262_nl = nl_MultLoop_acc_1262_nl[17:0];
  assign nl_MultLoop_acc_1375_nl = conv_s2u_20_21({(~ (data_rsci_idat[107:90])) ,
      2'b01}) + conv_s2u_19_21(MultLoop_acc_554_itm_23_5_1);
  assign MultLoop_acc_1375_nl = nl_MultLoop_acc_1375_nl[20:0];
  assign nl_MultLoop_acc_1263_nl = conv_s2u_19_20(readslicef_21_19_2((MultLoop_acc_1375_nl)))
      + ({(data_rsci_idat[107:90]) , 2'b01});
  assign MultLoop_acc_1263_nl = nl_MultLoop_acc_1263_nl[19:0];
  assign nl_MultLoop_acc_255_nl = conv_s2s_18_23(~ (data_rsci_idat[161:144])) + ({(data_rsci_idat[161:144])
      , 5'b00001});
  assign MultLoop_acc_255_nl = nl_MultLoop_acc_255_nl[22:0];
  assign nl_res_rsci_d_413_396  = (MultLoop_acc_553_nl) + conv_s2s_17_18(readslicef_22_17_5((MultLoop_acc_363_nl)))
      + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_1262_nl))) + conv_s2s_17_18(readslicef_20_17_3((MultLoop_acc_1263_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_255_nl)));
  assign nl_MultLoop_acc_1248_nl = (MultLoop_acc_901_itm_22_5[17:1]) + (~ (data_rsci_idat[52:36]));
  assign MultLoop_acc_1248_nl = nl_MultLoop_acc_1248_nl[16:0];
  assign nl_MultLoop_acc_903_nl = ({(data_rsci_idat[179:162]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_216_18_8
      , (~ (data_rsci_idat[169:162]))});
  assign MultLoop_acc_903_nl = nl_MultLoop_acc_903_nl[20:0];
  assign nl_MultLoop_acc_1250_nl = (~ (data_rsci_idat[179:162])) + conv_s2s_15_18(readslicef_21_15_6((MultLoop_acc_903_nl)));
  assign MultLoop_acc_1250_nl = nl_MultLoop_acc_1250_nl[17:0];
  assign nl_MultLoop_acc_1251_nl = conv_s2u_18_21(MultLoop_acc_1250_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[179:162])) , 2'b01});
  assign MultLoop_acc_1251_nl = nl_MultLoop_acc_1251_nl[20:0];
  assign nl_MultLoop_acc_911_nl = ({(MultLoop_acc_1248_nl) , (MultLoop_acc_901_itm_22_5[0])})
      + (readslicef_21_18_3((MultLoop_acc_1251_nl)));
  assign MultLoop_acc_911_nl = nl_MultLoop_acc_911_nl[17:0];
  assign nl_MultLoop_acc_111_nl = conv_s2u_15_18(data_rsci_idat[35:21]) - (data_rsci_idat[35:18]);
  assign MultLoop_acc_111_nl = nl_MultLoop_acc_111_nl[17:0];
  assign nl_MultLoop_acc_905_nl = conv_s2s_14_15(readslicef_18_14_4((MultLoop_acc_111_nl)))
      + 15'b000001110011101;
  assign MultLoop_acc_905_nl = nl_MultLoop_acc_905_nl[14:0];
  assign nl_MultLoop_acc_907_nl = MultLoop_acc_1348_itm_18_3 + conv_s2s_15_16(MultLoop_acc_905_nl);
  assign MultLoop_acc_907_nl = nl_MultLoop_acc_907_nl[15:0];
  assign nl_MultLoop_acc_1252_nl = (~ (data_rsci_idat[161:144])) + conv_s2s_16_18(MultLoop_acc_1374_itm_18_1[17:2]);
  assign MultLoop_acc_1252_nl = nl_MultLoop_acc_1252_nl[17:0];
  assign nl_MultLoop_acc_1253_nl = conv_s2u_18_20(MultLoop_acc_1252_nl) + ({(data_rsci_idat[161:144])
      , 2'b01});
  assign MultLoop_acc_1253_nl = nl_MultLoop_acc_1253_nl[19:0];
  assign nl_MultLoop_acc_910_nl = conv_s2s_16_18(MultLoop_acc_907_nl) + conv_s2s_17_18(readslicef_20_17_3((MultLoop_acc_1253_nl)));
  assign MultLoop_acc_910_nl = nl_MultLoop_acc_910_nl[17:0];
  assign nl_MultLoop_acc_913_nl = (MultLoop_acc_911_nl) + (MultLoop_acc_910_nl);
  assign MultLoop_acc_913_nl = nl_MultLoop_acc_913_nl[17:0];
  assign nl_MultLoop_acc_117_nl = conv_s2s_18_22(~ (data_rsci_idat[143:126])) + ({(data_rsci_idat[143:126])
      , 4'b0001});
  assign MultLoop_acc_117_nl = nl_MultLoop_acc_117_nl[21:0];
  assign nl_MultLoop_acc_891_nl = conv_s2s_18_19(data_rsci_idat[17:0]) + conv_s2s_17_19({MultLoop_acc_1254_cse_1
      , (data_rsci_idat[6:2])});
  assign MultLoop_acc_891_nl = nl_MultLoop_acc_891_nl[18:0];
  assign nl_MultLoop_acc_110_nl = conv_s2u_19_23(MultLoop_acc_891_nl) + ({(~ (data_rsci_idat[17:0]))
      , 5'b00000});
  assign MultLoop_acc_110_nl = nl_MultLoop_acc_110_nl[22:0];
  assign nl_MultLoop_acc_906_nl = conv_s2s_15_16(readslicef_22_15_7((MultLoop_acc_117_nl)))
      + conv_s2s_15_16(readslicef_23_15_8((MultLoop_acc_110_nl)));
  assign MultLoop_acc_906_nl = nl_MultLoop_acc_906_nl[15:0];
  assign nl_MultLoop_acc_908_nl = MultLoop_acc_302_itm_23_7 + conv_s2s_16_17(MultLoop_acc_906_nl);
  assign MultLoop_acc_908_nl = nl_MultLoop_acc_908_nl[16:0];
  assign nl_MultLoop_acc_896_nl = ({(data_rsci_idat[125:108]) , 3'b001}) + conv_s2s_18_21(MultLoop_acc_847_cse_1);
  assign MultLoop_acc_896_nl = nl_MultLoop_acc_896_nl[20:0];
  assign nl_MultLoop_acc_897_nl = ({(~ (data_rsci_idat[125:108])) , 5'b00000}) +
      conv_s2s_21_23(MultLoop_acc_896_nl);
  assign MultLoop_acc_897_nl = nl_MultLoop_acc_897_nl[22:0];
  assign nl_MultLoop_acc_324_nl = conv_s2u_23_25(MultLoop_acc_897_nl) + ({(data_rsci_idat[125:108])
      , 7'b0100000});
  assign MultLoop_acc_324_nl = nl_MultLoop_acc_324_nl[24:0];
  assign nl_MultLoop_acc_912_nl = conv_s2s_17_18(MultLoop_acc_908_nl) + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_324_nl)))
      + conv_s2s_17_18(MultLoop_acc_114_itm_19_3);
  assign MultLoop_acc_912_nl = nl_MultLoop_acc_912_nl[17:0];
  assign nl_res_rsci_d_179_162  = (MultLoop_acc_913_nl) + (MultLoop_acc_912_nl);
  assign nl_MultLoop_acc_1391_nl = conv_s2u_19_21(MultLoop_acc_1390_itm_22_4_1) +
      ({(data_rsci_idat[161:144]) , 3'b001});
  assign MultLoop_acc_1391_nl = nl_MultLoop_acc_1391_nl[20:0];
  assign nl_MultLoop_acc_567_nl = (~ (data_rsci_idat[179:162])) + conv_s2s_13_18(data_rsci_idat[179:167]);
  assign MultLoop_acc_567_nl = nl_MultLoop_acc_567_nl[17:0];
  assign nl_MultLoop_acc_568_nl = conv_s2s_20_21({(~ (data_rsci_idat[179:162])) ,
      2'b01}) + conv_s2s_18_21(MultLoop_acc_567_nl);
  assign MultLoop_acc_568_nl = nl_MultLoop_acc_568_nl[20:0];
  assign nl_MultLoop_acc_359_nl = conv_s2u_21_23(MultLoop_acc_568_nl) + ({(data_rsci_idat[179:162])
      , 5'b00100});
  assign MultLoop_acc_359_nl = nl_MultLoop_acc_359_nl[22:0];
  assign nl_MultLoop_acc_575_nl = (readslicef_21_18_3((MultLoop_acc_1391_nl))) +
      (readslicef_23_18_5((MultLoop_acc_359_nl)));
  assign MultLoop_acc_575_nl = nl_MultLoop_acc_575_nl[17:0];
  assign nl_MultLoop_acc_1371_nl = conv_s2u_17_19(MultLoop_acc_751_itm_18_2) + conv_s2u_18_19(data_rsci_idat[125:108]);
  assign MultLoop_acc_1371_nl = nl_MultLoop_acc_1371_nl[18:0];
  assign nl_MultLoop_acc_1372_nl = conv_s2u_19_20(MultLoop_acc_578_cse_1[21:3]) +
      ({(data_rsci_idat[89:72]) , 2'b01});
  assign MultLoop_acc_1372_nl = nl_MultLoop_acc_1372_nl[19:0];
  assign nl_MultLoop_acc_356_nl = conv_s2u_18_23(MultLoop_acc_557_cse_1) + ({(data_rsci_idat[35:18])
      , 5'b00001});
  assign MultLoop_acc_356_nl = nl_MultLoop_acc_356_nl[22:0];
  assign nl_MultLoop_acc_569_nl = conv_s2s_14_15(MultLoop_acc_237_itm_22_9) + 15'b000000111011001;
  assign MultLoop_acc_569_nl = nl_MultLoop_acc_569_nl[14:0];
  assign nl_MultLoop_acc_1370_nl = conv_s2u_19_20(MultLoop_acc_554_itm_23_5_1) +
      ({(data_rsci_idat[107:90]) , 2'b01});
  assign MultLoop_acc_1370_nl = nl_MultLoop_acc_1370_nl[19:0];
  assign nl_MultLoop_acc_574_nl = conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_1371_nl)))
      + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_1372_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_356_nl)))
      + conv_s2s_15_18(MultLoop_acc_569_nl) + conv_s2s_15_18(readslicef_20_15_5((MultLoop_acc_1370_nl)));
  assign MultLoop_acc_574_nl = nl_MultLoop_acc_574_nl[17:0];
  assign nl_MultLoop_acc_577_nl = (MultLoop_acc_575_nl) + (MultLoop_acc_574_nl);
  assign MultLoop_acc_577_nl = nl_MultLoop_acc_577_nl[17:0];
  assign nl_MultLoop_acc_240_nl = conv_s2s_27_28({(~ (data_rsci_idat[71:54])) , 9'b001000000})
      + conv_s2s_24_28({(~ (data_rsci_idat[71:54])) , 6'b000100}) + conv_s2s_20_28({(~
      (data_rsci_idat[71:54])) , 2'b01}) + conv_s2s_19_28({MultLoop_MultLoop_conc_228_18_9
      , (~ (data_rsci_idat[62:54]))});
  assign MultLoop_acc_240_nl = nl_MultLoop_acc_240_nl[27:0];
  assign nl_MultLoop_acc_558_nl = (~ (data_rsci_idat[143:126])) + conv_s2s_16_18(data_rsci_idat[143:128]);
  assign MultLoop_acc_558_nl = nl_MultLoop_acc_558_nl[17:0];
  assign nl_MultLoop_acc_559_nl = conv_s2s_21_22({(~ (data_rsci_idat[143:126])) ,
      3'b001}) + conv_s2s_18_22(MultLoop_acc_558_nl);
  assign MultLoop_acc_559_nl = nl_MultLoop_acc_559_nl[21:0];
  assign nl_MultLoop_acc_358_nl = conv_s2u_22_24(MultLoop_acc_559_nl) + ({(data_rsci_idat[143:126])
      , 6'b001000});
  assign MultLoop_acc_358_nl = nl_MultLoop_acc_358_nl[23:0];
  assign nl_MultLoop_acc_1373_nl = ({(data_rsci_idat[53:36]) , 3'b001}) + conv_s2u_19_21(MultLoop_acc_560_cse_1[21:3]);
  assign MultLoop_acc_1373_nl = nl_MultLoop_acc_1373_nl[20:0];
  assign nl_MultLoop_acc_1245_nl = conv_s2u_16_19(readslicef_21_16_5((MultLoop_acc_1373_nl)))
      + conv_s2u_18_19(data_rsci_idat[53:36]);
  assign MultLoop_acc_1245_nl = nl_MultLoop_acc_1245_nl[18:0];
  assign nl_res_rsci_d_395_378  = (MultLoop_acc_577_nl) + (readslicef_28_18_10((MultLoop_acc_240_nl)))
      + conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_358_nl))) + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_1245_nl)));
  assign nl_MultLoop_acc_1368_nl = ({(data_rsci_idat[125:108]) , 3'b001}) + conv_s2u_19_21(MultLoop_acc_1359_itm_20_2_1);
  assign MultLoop_acc_1368_nl = nl_MultLoop_acc_1368_nl[20:0];
  assign nl_MultLoop_acc_1237_nl = conv_s2u_16_19(readslicef_21_16_5((MultLoop_acc_1368_nl)))
      + conv_s2u_18_19(data_rsci_idat[125:108]);
  assign MultLoop_acc_1237_nl = nl_MultLoop_acc_1237_nl[18:0];
  assign nl_MultLoop_acc_880_nl = ({(data_rsci_idat[143:126]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[143:126]));
  assign MultLoop_acc_880_nl = nl_MultLoop_acc_880_nl[19:0];
  assign nl_MultLoop_acc_127_nl = conv_s2s_20_24(MultLoop_acc_880_nl) + conv_s2s_23_24({(data_rsci_idat[143:126])
      , 5'b00000});
  assign MultLoop_acc_127_nl = nl_MultLoop_acc_127_nl[23:0];
  assign nl_MultLoop_acc_887_nl = (readslicef_19_18_1((MultLoop_acc_1237_nl))) +
      (readslicef_24_18_6((MultLoop_acc_127_nl)));
  assign MultLoop_acc_887_nl = nl_MultLoop_acc_887_nl[17:0];
  assign nl_MultLoop_acc_881_nl = ({(data_rsci_idat[161:144]) , 4'b0001}) + conv_s2s_18_22(~
      (data_rsci_idat[161:144]));
  assign MultLoop_acc_881_nl = nl_MultLoop_acc_881_nl[21:0];
  assign nl_MultLoop_acc_1238_nl = conv_s2u_14_19(readslicef_22_14_8((MultLoop_acc_881_nl)))
      + conv_s2u_18_19(data_rsci_idat[161:144]);
  assign MultLoop_acc_1238_nl = nl_MultLoop_acc_1238_nl[18:0];
  assign nl_MultLoop_acc_867_nl = conv_s2s_18_19(data_rsci_idat[17:0]) + conv_s2s_17_19({MultLoop_acc_1239_cse_1
      , (data_rsci_idat[4:2])});
  assign MultLoop_acc_867_nl = nl_MultLoop_acc_867_nl[18:0];
  assign nl_MultLoop_acc_120_nl = conv_s2u_19_21(MultLoop_acc_867_nl) + ({(~ (data_rsci_idat[17:0]))
      , 3'b000});
  assign MultLoop_acc_120_nl = nl_MultLoop_acc_120_nl[20:0];
  assign nl_MultLoop_101_MultLoop_acc_3_nl = (readslicef_21_15_6((MultLoop_acc_120_nl)))
      + 15'b000000110100111;
  assign MultLoop_101_MultLoop_acc_3_nl = nl_MultLoop_101_MultLoop_acc_3_nl[14:0];
  assign nl_MultLoop_acc_124_nl = conv_s2u_16_18(data_rsci_idat[89:74]) - (data_rsci_idat[89:72]);
  assign MultLoop_acc_124_nl = nl_MultLoop_acc_124_nl[17:0];
  assign nl_MultLoop_acc_884_nl = conv_s2s_16_17(MultLoop_acc_620_itm_18_3) + conv_s2s_15_17(MultLoop_101_MultLoop_acc_3_nl)
      + conv_s2s_13_17(MultLoop_acc_123_itm_21_6[15:3]) + conv_s2s_12_17(readslicef_18_12_6((MultLoop_acc_124_nl)));
  assign MultLoop_acc_884_nl = nl_MultLoop_acc_884_nl[16:0];
  assign nl_MultLoop_acc_886_nl = (readslicef_19_18_1((MultLoop_acc_1238_nl))) +
      conv_s2s_17_18(MultLoop_acc_884_nl);
  assign MultLoop_acc_886_nl = nl_MultLoop_acc_886_nl[17:0];
  assign nl_MultLoop_acc_889_nl = (MultLoop_acc_887_nl) + (MultLoop_acc_886_nl);
  assign MultLoop_acc_889_nl = nl_MultLoop_acc_889_nl[17:0];
  assign nl_MultLoop_acc_1240_nl =  -conv_s2s_9_10(data_rsci_idat[179:171]);
  assign MultLoop_acc_1240_nl = nl_MultLoop_acc_1240_nl[9:0];
  assign nl_MultLoop_acc_869_nl = ({(data_rsci_idat[179:162]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_1240_nl)
      , (~ (data_rsci_idat[170:162]))});
  assign MultLoop_acc_869_nl = nl_MultLoop_acc_869_nl[19:0];
  assign nl_MultLoop_acc_870_nl = ({(~ (data_rsci_idat[179:162])) , 4'b0000}) + conv_s2s_20_22(MultLoop_acc_869_nl);
  assign MultLoop_acc_870_nl = nl_MultLoop_acc_870_nl[21:0];
  assign nl_MultLoop_acc_871_nl = ({(data_rsci_idat[179:162]) , 6'b010000}) + conv_s2s_22_24(MultLoop_acc_870_nl);
  assign MultLoop_acc_871_nl = nl_MultLoop_acc_871_nl[23:0];
  assign nl_MultLoop_acc_1241_nl = conv_s2u_15_18(readslicef_24_15_9((MultLoop_acc_871_nl)))
      + (~ (data_rsci_idat[179:162]));
  assign MultLoop_acc_1241_nl = nl_MultLoop_acc_1241_nl[17:0];
  assign nl_MultLoop_acc_874_nl = ({(data_rsci_idat[53:36]) , 6'b010000}) + conv_s2s_22_24({(~
      (data_rsci_idat[53:36])) , 4'b0001}) + conv_s2s_19_24({MultLoop_MultLoop_conc_218_18_8
      , (~ (data_rsci_idat[43:36]))});
  assign MultLoop_acc_874_nl = nl_MultLoop_acc_874_nl[23:0];
  assign nl_MultLoop_acc_1243_nl = conv_s2u_16_18(readslicef_24_16_8((MultLoop_acc_874_nl)))
      + (~ (data_rsci_idat[53:36]));
  assign MultLoop_acc_1243_nl = nl_MultLoop_acc_1243_nl[17:0];
  assign nl_MultLoop_acc_885_nl = conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_1241_nl)))
      + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_1243_nl)));
  assign MultLoop_acc_885_nl = nl_MultLoop_acc_885_nl[17:0];
  assign nl_MultLoop_acc_1369_nl = conv_s2u_18_19(data_rsci_idat[35:18]) + conv_s2u_17_19(MultLoop_acc_875_cse_1[18:2]);
  assign MultLoop_acc_1369_nl = nl_MultLoop_acc_1369_nl[18:0];
  assign nl_MultLoop_acc_1244_nl = conv_s2u_14_19(readslicef_19_14_5((MultLoop_acc_1369_nl)))
      + conv_s2u_18_19(data_rsci_idat[35:18]);
  assign MultLoop_acc_1244_nl = nl_MultLoop_acc_1244_nl[18:0];
  assign nl_MultLoop_acc_888_nl = (MultLoop_acc_885_nl) + (readslicef_19_18_1((MultLoop_acc_1244_nl)));
  assign MultLoop_acc_888_nl = nl_MultLoop_acc_888_nl[17:0];
  assign nl_res_rsci_d_197_180  = (MultLoop_acc_889_nl) + (MultLoop_acc_888_nl);
  assign nl_MultLoop_acc_587_nl = ({(data_rsci_idat[125:108]) , 7'b0010000}) + conv_s2s_22_25({(~
      (data_rsci_idat[125:108])) , 4'b0100}) + conv_s2s_20_25({(~ (data_rsci_idat[125:108]))
      , 2'b01}) + conv_s2s_19_25({MultLoop_MultLoop_conc_222_18_9 , (~ (data_rsci_idat[116:108]))});
  assign MultLoop_acc_587_nl = nl_MultLoop_acc_587_nl[24:0];
  assign nl_MultLoop_acc_1233_nl = conv_s2u_16_18(readslicef_25_16_9((MultLoop_acc_587_nl)))
      + (~ (data_rsci_idat[125:108]));
  assign MultLoop_acc_1233_nl = nl_MultLoop_acc_1233_nl[17:0];
  assign nl_MultLoop_acc_591_nl = ({(data_rsci_idat[143:126]) , 7'b0100000}) + conv_s2s_23_25({(~
      (data_rsci_idat[143:126])) , 5'b00100}) + conv_s2s_20_25({(~ (data_rsci_idat[143:126]))
      , 2'b01}) + conv_s2s_19_25({Result_Result_conc_48_18_9 , (~ (data_rsci_idat[134:126]))});
  assign MultLoop_acc_591_nl = nl_MultLoop_acc_591_nl[24:0];
  assign nl_MultLoop_acc_1235_nl = conv_s2u_16_18(readslicef_25_16_9((MultLoop_acc_591_nl)))
      + (~ (data_rsci_idat[143:126]));
  assign MultLoop_acc_1235_nl = nl_MultLoop_acc_1235_nl[17:0];
  assign nl_MultLoop_acc_1236_nl =  -conv_s2s_13_14(data_rsci_idat[35:23]);
  assign MultLoop_acc_1236_nl = nl_MultLoop_acc_1236_nl[13:0];
  assign nl_MultLoop_acc_229_nl = conv_s2s_23_24({(~ (data_rsci_idat[35:18])) , 5'b01000})
      + conv_s2s_21_24({(~ (data_rsci_idat[35:18])) , 3'b001}) + conv_s2s_19_24({(MultLoop_acc_1236_nl)
      , (~ (data_rsci_idat[22:18]))});
  assign MultLoop_acc_229_nl = nl_MultLoop_acc_229_nl[23:0];
  assign nl_MultLoop_acc_595_nl = (readslicef_24_16_8((MultLoop_acc_229_nl))) + 16'b0000000001110101;
  assign MultLoop_acc_595_nl = nl_MultLoop_acc_595_nl[15:0];
  assign nl_MultLoop_acc_1407_nl = conv_s2u_17_19(MultLoop_acc_594_itm_18_2_1) +
      conv_s2u_18_19(data_rsci_idat[17:0]);
  assign MultLoop_acc_1407_nl = nl_MultLoop_acc_1407_nl[18:0];
  assign nl_MultLoop_202_MultLoop_acc_3_nl = conv_s2s_16_17(MultLoop_acc_595_nl)
      + (readslicef_19_17_2((MultLoop_acc_1407_nl)));
  assign MultLoop_202_MultLoop_acc_3_nl = nl_MultLoop_202_MultLoop_acc_3_nl[16:0];
  assign nl_MultLoop_acc_603_nl = conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_1233_nl)))
      + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_1235_nl))) + conv_s2s_17_18(MultLoop_202_MultLoop_acc_3_nl)
      + conv_s2s_17_18(MultLoop_acc_353_itm_22_6);
  assign MultLoop_acc_603_nl = nl_MultLoop_acc_603_nl[17:0];
  assign nl_MultLoop_acc_1367_nl = conv_s2u_18_19(data_rsci_idat[53:36]) + conv_s2u_16_19(MultLoop_acc_596_itm_20_5);
  assign MultLoop_acc_1367_nl = nl_MultLoop_acc_1367_nl[18:0];
  assign nl_MultLoop_acc_1231_nl = conv_s2u_17_19(readslicef_19_17_2((MultLoop_acc_1367_nl)))
      + conv_s2u_18_19(data_rsci_idat[53:36]);
  assign MultLoop_acc_1231_nl = nl_MultLoop_acc_1231_nl[18:0];
  assign nl_MultLoop_acc_579_nl = conv_s2s_23_24({(~ (data_rsci_idat[89:72])) , 5'b01000})
      + conv_s2s_22_24(MultLoop_acc_578_cse_1);
  assign MultLoop_acc_579_nl = nl_MultLoop_acc_579_nl[23:0];
  assign nl_MultLoop_acc_232_nl = conv_s2s_24_26(MultLoop_acc_579_nl) + ({(data_rsci_idat[89:72])
      , 8'b00100000});
  assign MultLoop_acc_232_nl = nl_MultLoop_acc_232_nl[25:0];
  assign nl_MultLoop_acc_598_nl = conv_s2s_16_17(readslicef_26_16_10((MultLoop_acc_232_nl)))
      + conv_s2s_15_17(data_rsci_idat[107:93]);
  assign MultLoop_acc_598_nl = nl_MultLoop_acc_598_nl[16:0];
  assign nl_MultLoop_acc_602_nl = (readslicef_19_18_1((MultLoop_acc_1231_nl))) +
      conv_s2s_17_18(MultLoop_acc_598_nl);
  assign MultLoop_acc_602_nl = nl_MultLoop_acc_602_nl[17:0];
  assign nl_MultLoop_acc_1409_nl = conv_s2u_15_19(MultLoop_acc_1401_itm_20_5[15:1])
      + conv_s2u_18_19(data_rsci_idat[161:144]);
  assign MultLoop_acc_1409_nl = nl_MultLoop_acc_1409_nl[18:0];
  assign nl_MultLoop_acc_1389_nl = conv_s2u_18_21(MultLoop_asn_361) + ({(data_rsci_idat[179:162])
      , 3'b001});
  assign MultLoop_acc_1389_nl = nl_MultLoop_acc_1389_nl[20:0];
  assign nl_res_rsci_d_377_360  = (MultLoop_acc_603_nl) + (MultLoop_acc_602_nl) +
      conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_1409_nl))) + conv_s2s_17_18(readslicef_21_17_4((MultLoop_acc_1389_nl)));
  assign nl_MultLoop_acc_1222_nl = conv_s2s_12_13(data_rsci_idat[89:78]) + 13'b0000000000001;
  assign MultLoop_acc_1222_nl = nl_MultLoop_acc_1222_nl[12:0];
  assign nl_MultLoop_acc_836_nl = ({(~ (data_rsci_idat[89:72])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[89:72])
      + conv_s2s_17_20({(MultLoop_acc_1222_nl) , (data_rsci_idat[77:74])});
  assign MultLoop_acc_836_nl = nl_MultLoop_acc_836_nl[19:0];
  assign nl_MultLoop_acc_327_nl = conv_s2u_20_23(MultLoop_acc_836_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[89:72])) , 4'b0100});
  assign MultLoop_acc_327_nl = nl_MultLoop_acc_327_nl[22:0];
  assign nl_MultLoop_acc_837_nl = (~ (data_rsci_idat[107:90])) + conv_s2s_14_18(data_rsci_idat[107:94]);
  assign MultLoop_acc_837_nl = nl_MultLoop_acc_837_nl[17:0];
  assign nl_MultLoop_acc_838_nl = ({(data_rsci_idat[107:90]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_837_nl);
  assign MultLoop_acc_838_nl = nl_MultLoop_acc_838_nl[19:0];
  assign nl_MultLoop_acc_328_nl = conv_s2u_20_23(MultLoop_acc_838_nl) + conv_s2u_22_23({(data_rsci_idat[107:90])
      , 4'b0000});
  assign MultLoop_acc_328_nl = nl_MultLoop_acc_328_nl[22:0];
  assign nl_MultLoop_acc_858_nl = conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_327_nl)))
      + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_328_nl)));
  assign MultLoop_acc_858_nl = nl_MultLoop_acc_858_nl[17:0];
  assign nl_MultLoop_acc_1366_nl = conv_s2u_23_24({(~ (data_rsci_idat[35:18])) ,
      5'b00001}) + conv_s2u_19_24(MultLoop_acc_839_cse_1[21:3]);
  assign MultLoop_acc_1366_nl = nl_MultLoop_acc_1366_nl[23:0];
  assign nl_MultLoop_acc_1223_nl = conv_s2u_19_20(readslicef_24_19_5((MultLoop_acc_1366_nl)))
      + ({(data_rsci_idat[35:18]) , 2'b01});
  assign MultLoop_acc_1223_nl = nl_MultLoop_acc_1223_nl[19:0];
  assign nl_MultLoop_acc_862_nl = (MultLoop_acc_858_nl) + (readslicef_20_18_2((MultLoop_acc_1223_nl)));
  assign MultLoop_acc_862_nl = nl_MultLoop_acc_862_nl[17:0];
  assign nl_MultLoop_acc_843_nl = ({(data_rsci_idat[53:36]) , 3'b001}) + conv_s2s_18_21(MultLoop_acc_642_cse_1);
  assign MultLoop_acc_843_nl = nl_MultLoop_acc_843_nl[20:0];
  assign nl_MultLoop_acc_133_nl = conv_s2u_21_23(MultLoop_acc_843_nl) + ({(~ (data_rsci_idat[53:36]))
      , 5'b00000});
  assign MultLoop_acc_133_nl = nl_MultLoop_acc_133_nl[22:0];
  assign nl_MultLoop_acc_845_nl = ({(data_rsci_idat[71:54]) , 2'b01}) + conv_s2s_19_20({Result_Result_conc_64_18_8
      , (~ (data_rsci_idat[61:54]))});
  assign MultLoop_acc_845_nl = nl_MultLoop_acc_845_nl[19:0];
  assign nl_MultLoop_acc_846_nl = ({(~ (data_rsci_idat[71:54])) , 4'b0000}) + conv_s2s_20_22(MultLoop_acc_845_nl);
  assign MultLoop_acc_846_nl = nl_MultLoop_acc_846_nl[21:0];
  assign nl_MultLoop_acc_134_nl = conv_s2s_22_27(MultLoop_acc_846_nl) + conv_s2s_26_27({(~
      (data_rsci_idat[71:54])) , 8'b00010000});
  assign MultLoop_acc_134_nl = nl_MultLoop_acc_134_nl[26:0];
  assign nl_MultLoop_acc_861_nl = (readslicef_23_18_5((MultLoop_acc_133_nl))) + (readslicef_27_18_9((MultLoop_acc_134_nl)));
  assign MultLoop_acc_861_nl = nl_MultLoop_acc_861_nl[17:0];
  assign nl_MultLoop_acc_864_nl = (MultLoop_acc_862_nl) + (MultLoop_acc_861_nl);
  assign MultLoop_acc_864_nl = nl_MultLoop_acc_864_nl[17:0];
  assign nl_MultLoop_acc_849_nl = ({(data_rsci_idat[125:108]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[125:108])) , 2'b01}) + conv_s2s_18_22(MultLoop_acc_847_cse_1);
  assign MultLoop_acc_849_nl = nl_MultLoop_acc_849_nl[21:0];
  assign nl_MultLoop_acc_329_nl = conv_s2u_22_25(MultLoop_acc_849_nl) + conv_s2u_24_25({(data_rsci_idat[125:108])
      , 6'b000000});
  assign MultLoop_acc_329_nl = nl_MultLoop_acc_329_nl[24:0];
  assign nl_MultLoop_acc_853_nl = conv_s2s_26_27({(~ (data_rsci_idat[161:144])) ,
      8'b00100000}) + conv_s2s_23_27({(~ (data_rsci_idat[161:144])) , 5'b00100})
      + conv_s2s_20_27({(~ (data_rsci_idat[161:144])) , 2'b01}) + conv_s2s_19_27({Result_Result_conc_52_18_10
      , (~ (data_rsci_idat[153:144]))});
  assign MultLoop_acc_853_nl = nl_MultLoop_acc_853_nl[26:0];
  assign nl_MultLoop_acc_1227_nl = conv_s2u_19_20(readslicef_27_19_8((MultLoop_acc_853_nl)))
      + ({(~ (data_rsci_idat[161:144])) , 2'b01});
  assign MultLoop_acc_1227_nl = nl_MultLoop_acc_1227_nl[19:0];
  assign nl_MultLoop_acc_860_nl = (readslicef_25_18_7((MultLoop_acc_329_nl))) + (readslicef_20_18_2((MultLoop_acc_1227_nl)));
  assign MultLoop_acc_860_nl = nl_MultLoop_acc_860_nl[17:0];
  assign nl_MultLoop_acc_1228_nl =  -conv_s2s_11_12(data_rsci_idat[179:169]);
  assign MultLoop_acc_1228_nl = nl_MultLoop_acc_1228_nl[11:0];
  assign nl_MultLoop_acc_855_nl = conv_s2s_21_22({(~ (data_rsci_idat[179:162])) ,
      3'b001}) + conv_s2s_19_22({(MultLoop_acc_1228_nl) , (~ (data_rsci_idat[168:162]))});
  assign MultLoop_acc_855_nl = nl_MultLoop_acc_855_nl[21:0];
  assign nl_MultLoop_acc_140_nl = conv_s2s_22_25(MultLoop_acc_855_nl) + ({(~ (data_rsci_idat[179:162]))
      , 7'b0001000});
  assign MultLoop_acc_140_nl = nl_MultLoop_acc_140_nl[24:0];
  assign nl_MultLoop_acc_832_nl = (~ (data_rsci_idat[143:126])) + conv_s2s_15_18(data_rsci_idat[143:129]);
  assign MultLoop_acc_832_nl = nl_MultLoop_acc_832_nl[17:0];
  assign nl_MultLoop_acc_833_nl = conv_s2s_21_22({(~ (data_rsci_idat[143:126])) ,
      3'b001}) + conv_s2s_18_22(MultLoop_acc_832_nl);
  assign MultLoop_acc_833_nl = nl_MultLoop_acc_833_nl[21:0];
  assign nl_MultLoop_acc_330_nl = conv_s2u_22_23(MultLoop_acc_833_nl) + ({(data_rsci_idat[143:126])
      , 5'b01000});
  assign MultLoop_acc_330_nl = nl_MultLoop_acc_330_nl[22:0];
  assign nl_MultLoop_acc_1230_nl = (MultLoop_acc_130_itm_20_10[10:1]) + 10'b0010010101;
  assign MultLoop_acc_1230_nl = nl_MultLoop_acc_1230_nl[9:0];
  assign nl_MultLoop_acc_859_nl = (readslicef_25_18_7((MultLoop_acc_140_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_330_nl)))
      + conv_s2s_11_18({(MultLoop_acc_1230_nl) , (MultLoop_acc_130_itm_20_10[0])});
  assign MultLoop_acc_859_nl = nl_MultLoop_acc_859_nl[17:0];
  assign nl_MultLoop_acc_863_nl = (MultLoop_acc_860_nl) + (MultLoop_acc_859_nl);
  assign MultLoop_acc_863_nl = nl_MultLoop_acc_863_nl[17:0];
  assign nl_res_rsci_d_215_198  = (MultLoop_acc_864_nl) + (MultLoop_acc_863_nl);
  assign nl_MultLoop_acc_1363_nl = conv_s2u_16_19(MultLoop_acc_620_itm_18_3) + conv_s2u_18_19(data_rsci_idat[107:90]);
  assign MultLoop_acc_1363_nl = nl_MultLoop_acc_1363_nl[18:0];
  assign nl_MultLoop_acc_622_nl = ({(data_rsci_idat[125:108]) , 4'b0001}) + conv_s2s_18_22(MultLoop_acc_621_cse_1);
  assign MultLoop_acc_622_nl = nl_MultLoop_acc_622_nl[21:0];
  assign nl_MultLoop_acc_352_nl = conv_s2u_22_25(MultLoop_acc_622_nl) + conv_s2u_24_25({(data_rsci_idat[125:108])
      , 6'b000000});
  assign MultLoop_acc_352_nl = nl_MultLoop_acc_352_nl[24:0];
  assign nl_MultLoop_acc_629_nl = (readslicef_19_18_1((MultLoop_acc_1363_nl))) +
      (readslicef_25_18_7((MultLoop_acc_352_nl)));
  assign MultLoop_acc_629_nl = nl_MultLoop_acc_629_nl[17:0];
  assign nl_MultLoop_acc_1364_nl = conv_s2u_16_19(MultLoop_acc_623_cse_1[20:5]) +
      conv_s2u_18_19(data_rsci_idat[143:126]);
  assign MultLoop_acc_1364_nl = nl_MultLoop_acc_1364_nl[18:0];
  assign nl_MultLoop_acc_618_nl = ({(data_rsci_idat[71:54]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_202_18_7
      , (~ (data_rsci_idat[60:54]))});
  assign MultLoop_acc_618_nl = nl_MultLoop_acc_618_nl[19:0];
  assign nl_MultLoop_acc_619_nl = ({(~ (data_rsci_idat[71:54])) , 5'b00000}) + conv_s2s_20_23(MultLoop_acc_618_nl);
  assign MultLoop_acc_619_nl = nl_MultLoop_acc_619_nl[22:0];
  assign nl_MultLoop_acc_220_nl = conv_s2s_23_26(MultLoop_acc_619_nl) + conv_s2s_25_26({(~
      (data_rsci_idat[71:54])) , 7'b0100000});
  assign MultLoop_acc_220_nl = nl_MultLoop_acc_220_nl[25:0];
  assign nl_MultLoop_acc_605_nl = conv_s2s_24_25({(~ (data_rsci_idat[89:72])) , 6'b000001})
      + conv_s2s_18_25(~ (data_rsci_idat[89:72]));
  assign MultLoop_acc_605_nl = nl_MultLoop_acc_605_nl[24:0];
  assign nl_MultLoop_acc_221_nl = conv_s2s_25_26(MultLoop_acc_605_nl) + ({(data_rsci_idat[89:72])
      , 8'b01000000});
  assign MultLoop_acc_221_nl = nl_MultLoop_acc_221_nl[25:0];
  assign nl_MultLoop_acc_625_nl = (readslicef_26_17_9((MultLoop_acc_220_nl))) + conv_s2s_16_17(readslicef_26_16_10((MultLoop_acc_221_nl)));
  assign MultLoop_acc_625_nl = nl_MultLoop_acc_625_nl[16:0];
  assign nl_MultLoop_acc_628_nl = (readslicef_19_18_1((MultLoop_acc_1364_nl))) +
      conv_s2s_17_18(MultLoop_acc_625_nl);
  assign MultLoop_acc_628_nl = nl_MultLoop_acc_628_nl[17:0];
  assign nl_MultLoop_acc_631_nl = (MultLoop_acc_629_nl) + (MultLoop_acc_628_nl);
  assign MultLoop_acc_631_nl = nl_MultLoop_acc_631_nl[17:0];
  assign nl_MultLoop_acc_225_nl = conv_s2s_24_25({(~ (data_rsci_idat[161:144])) ,
      6'b000100}) + conv_s2s_20_25({(~ (data_rsci_idat[161:144])) , 2'b01}) + conv_s2s_19_25({MultLoop_MultLoop_conc_212_18_6
      , (~ (data_rsci_idat[149:144]))});
  assign MultLoop_acc_225_nl = nl_MultLoop_acc_225_nl[24:0];
  assign nl_MultLoop_acc_1365_nl = conv_s2u_15_19(MultLoop_acc_731_itm_18_4) + conv_s2u_18_19(data_rsci_idat[17:0]);
  assign MultLoop_acc_1365_nl = nl_MultLoop_acc_1365_nl[18:0];
  assign nl_MultLoop_191_MultLoop_acc_3_nl = (readslicef_19_16_3((MultLoop_acc_1365_nl)))
      + 16'b1111111101010111;
  assign MultLoop_191_MultLoop_acc_3_nl = nl_MultLoop_191_MultLoop_acc_3_nl[15:0];
  assign nl_MultLoop_acc_608_nl = ({(data_rsci_idat[35:18]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[35:18])) , 2'b01}) + conv_s2s_18_22(~ (data_rsci_idat[35:18]));
  assign MultLoop_acc_608_nl = nl_MultLoop_acc_608_nl[21:0];
  assign nl_MultLoop_acc_1217_nl = (~ (data_rsci_idat[35:18])) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_608_nl)));
  assign MultLoop_acc_1217_nl = nl_MultLoop_acc_1217_nl[17:0];
  assign nl_MultLoop_acc_1218_nl = conv_s2u_18_20(MultLoop_acc_1217_nl) + ({(data_rsci_idat[35:18])
      , 2'b01});
  assign MultLoop_acc_1218_nl = nl_MultLoop_acc_1218_nl[19:0];
  assign nl_MultLoop_acc_1220_nl =  -conv_s2s_12_13(data_rsci_idat[179:168]);
  assign MultLoop_acc_1220_nl = nl_MultLoop_acc_1220_nl[12:0];
  assign nl_MultLoop_acc_613_nl = ({(data_rsci_idat[179:162]) , 4'b0001}) + conv_s2s_19_22({(MultLoop_acc_1220_nl)
      , (~ (data_rsci_idat[167:162]))});
  assign MultLoop_acc_613_nl = nl_MultLoop_acc_613_nl[21:0];
  assign nl_MultLoop_acc_1221_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_613_nl)))
      + (~ (data_rsci_idat[179:162]));
  assign MultLoop_acc_1221_nl = nl_MultLoop_acc_1221_nl[17:0];
  assign nl_MultLoop_acc_614_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_16_18(data_rsci_idat[53:38]);
  assign MultLoop_acc_614_nl = nl_MultLoop_acc_614_nl[17:0];
  assign nl_MultLoop_acc_615_nl = ({(data_rsci_idat[53:36]) , 3'b001}) + conv_s2s_18_21(MultLoop_acc_614_nl);
  assign MultLoop_acc_615_nl = nl_MultLoop_acc_615_nl[20:0];
  assign nl_MultLoop_acc_616_nl = ({(~ (data_rsci_idat[53:36])) , 5'b00000}) + conv_s2s_21_23(MultLoop_acc_615_nl);
  assign MultLoop_acc_616_nl = nl_MultLoop_acc_616_nl[22:0];
  assign nl_MultLoop_acc_350_nl = conv_s2u_23_25(MultLoop_acc_616_nl) + ({(data_rsci_idat[53:36])
      , 7'b0100000});
  assign MultLoop_acc_350_nl = nl_MultLoop_acc_350_nl[24:0];
  assign nl_res_rsci_d_359_342  = (MultLoop_acc_631_nl) + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_225_nl)))
      + conv_s2s_16_18(MultLoop_191_MultLoop_acc_3_nl) + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_1218_nl)))
      + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_1221_nl))) + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_350_nl)));
  assign nl_MultLoop_acc_1362_nl = conv_s2u_19_20(MultLoop_acc_660_itm_22_4_1) +
      ({(data_rsci_idat[89:72]) , 2'b01});
  assign MultLoop_acc_1362_nl = nl_MultLoop_acc_1362_nl[19:0];
  assign nl_MultLoop_acc_813_nl = ({(~ (data_rsci_idat[35:18])) , 2'b00}) + conv_s2s_19_20(MultLoop_acc_812_cse_1);
  assign MultLoop_acc_813_nl = nl_MultLoop_acc_813_nl[19:0];
  assign nl_MultLoop_acc_331_nl = conv_s2u_20_22(MultLoop_acc_813_nl) + ({(data_rsci_idat[35:18])
      , 4'b0100});
  assign MultLoop_acc_331_nl = nl_MultLoop_acc_331_nl[21:0];
  assign nl_MultLoop_acc_1212_nl = conv_s2s_13_14(data_rsci_idat[107:95]) + 14'b00000000000001;
  assign MultLoop_acc_1212_nl = nl_MultLoop_acc_1212_nl[13:0];
  assign nl_MultLoop_acc_804_nl = (~ (data_rsci_idat[107:90])) + conv_s2s_17_18({(MultLoop_acc_1212_nl)
      , (data_rsci_idat[94:92])});
  assign MultLoop_acc_804_nl = nl_MultLoop_acc_804_nl[17:0];
  assign nl_MultLoop_acc_332_nl = conv_s2u_18_22(MultLoop_acc_804_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[107:90])) , 3'b001});
  assign MultLoop_acc_332_nl = nl_MultLoop_acc_332_nl[21:0];
  assign nl_MultLoop_acc_822_nl = (readslicef_22_14_8((MultLoop_acc_332_nl))) + 14'b00000010111111;
  assign MultLoop_acc_822_nl = nl_MultLoop_acc_822_nl[13:0];
  assign nl_MultLoop_acc_1210_nl = conv_s2s_11_12(data_rsci_idat[179:169]) + 12'b000000000001;
  assign MultLoop_acc_1210_nl = nl_MultLoop_acc_1210_nl[11:0];
  assign nl_MultLoop_acc_807_nl = (~ (data_rsci_idat[179:162])) + conv_s2s_16_18({(MultLoop_acc_1210_nl)
      , (data_rsci_idat[168:165])});
  assign MultLoop_acc_807_nl = nl_MultLoop_acc_807_nl[17:0];
  assign nl_MultLoop_acc_334_nl = conv_s2u_18_23(MultLoop_acc_807_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[179:162])) , 4'b0001});
  assign MultLoop_acc_334_nl = nl_MultLoop_acc_334_nl[22:0];
  assign nl_MultLoop_acc_1360_nl = conv_s2u_14_19(MultLoop_acc_805_cse_1[19:6]) +
      conv_s2u_18_19(data_rsci_idat[17:0]);
  assign MultLoop_acc_1360_nl = nl_MultLoop_acc_1360_nl[18:0];
  assign nl_MultLoop_acc_1361_nl = conv_s2u_19_22(MultLoop_acc_1359_itm_20_2_1) +
      ({(data_rsci_idat[125:108]) , 4'b0001});
  assign MultLoop_acc_1361_nl = nl_MultLoop_acc_1361_nl[21:0];
  assign nl_MultLoop_acc_811_nl = conv_s2s_18_19(data_rsci_idat[53:36]) + conv_s2s_14_19({Result_Result_conc_50_13_2
      , (data_rsci_idat[42:41])});
  assign MultLoop_acc_811_nl = nl_MultLoop_acc_811_nl[18:0];
  assign nl_MultLoop_acc_143_nl = conv_s2u_19_20(MultLoop_acc_811_nl) + ({(~ (data_rsci_idat[53:36]))
      , 2'b00});
  assign MultLoop_acc_143_nl = nl_MultLoop_acc_143_nl[19:0];
  assign nl_MultLoop_acc_830_nl = conv_s2s_17_18(readslicef_20_17_3((MultLoop_acc_1362_nl)))
      + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_331_nl))) + conv_s2s_14_18(MultLoop_acc_822_nl)
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_334_nl))) + conv_s2s_15_18(readslicef_19_15_4((MultLoop_acc_1360_nl)))
      + conv_s2s_14_18(MultLoop_acc_74_itm_17_1[16:3]) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1361_nl)))
      + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_143_nl)));
  assign MultLoop_acc_830_nl = nl_MultLoop_acc_830_nl[17:0];
  assign nl_MultLoop_acc_816_nl = (~ (data_rsci_idat[71:54])) + conv_s2s_17_18({MultLoop_acc_1213_cse_1
      , (data_rsci_idat[63:56])});
  assign MultLoop_acc_816_nl = nl_MultLoop_acc_816_nl[17:0];
  assign nl_MultLoop_acc_818_nl = ({(data_rsci_idat[71:54]) , 6'b000100}) + conv_s2s_20_24({(~
      (data_rsci_idat[71:54])) , 2'b01}) + conv_s2s_18_24(MultLoop_acc_816_nl);
  assign MultLoop_acc_818_nl = nl_MultLoop_acc_818_nl[23:0];
  assign nl_MultLoop_acc_1214_nl = conv_s2u_16_18(readslicef_24_16_8((MultLoop_acc_818_nl)))
      + (~ (data_rsci_idat[71:54]));
  assign MultLoop_acc_1214_nl = nl_MultLoop_acc_1214_nl[17:0];
  assign nl_MultLoop_acc_1408_nl = conv_s2u_18_19(data_rsci_idat[161:144]) + conv_s2u_16_19(MultLoop_acc_1401_itm_20_5);
  assign MultLoop_acc_1408_nl = nl_MultLoop_acc_1408_nl[18:0];
  assign nl_MultLoop_acc_1215_nl = conv_s2u_16_18(readslicef_19_16_3((MultLoop_acc_1408_nl)))
      + (data_rsci_idat[161:144]);
  assign MultLoop_acc_1215_nl = nl_MultLoop_acc_1215_nl[17:0];
  assign nl_MultLoop_acc_829_nl = (MultLoop_acc_1214_nl) + (MultLoop_acc_1215_nl);
  assign MultLoop_acc_829_nl = nl_MultLoop_acc_829_nl[17:0];
  assign nl_res_rsci_d_233_216  = (MultLoop_acc_830_nl) + (MultLoop_acc_829_nl);
  assign nl_MultLoop_acc_643_nl = ({(data_rsci_idat[53:36]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_642_cse_1);
  assign MultLoop_acc_643_nl = nl_MultLoop_acc_643_nl[19:0];
  assign nl_MultLoop_acc_208_nl = conv_s2u_20_23(MultLoop_acc_643_nl) + ({(~ (data_rsci_idat[53:36]))
      , 5'b00000});
  assign MultLoop_acc_208_nl = nl_MultLoop_acc_208_nl[22:0];
  assign nl_MultLoop_acc_209_nl = conv_s2s_27_28({(~ (data_rsci_idat[71:54])) , 9'b000010000})
      + conv_s2s_22_28({(~ (data_rsci_idat[71:54])) , 4'b0001}) + conv_s2s_19_28({MultLoop_MultLoop_conc_228_18_9
      , (~ (data_rsci_idat[62:54]))});
  assign MultLoop_acc_209_nl = nl_MultLoop_acc_209_nl[27:0];
  assign nl_MultLoop_acc_657_nl = (readslicef_23_18_5((MultLoop_acc_208_nl))) + (readslicef_28_18_10((MultLoop_acc_209_nl)));
  assign MultLoop_acc_657_nl = nl_MultLoop_acc_657_nl[17:0];
  assign nl_MultLoop_acc_1205_nl = conv_s2s_9_10(data_rsci_idat[89:81]) + 10'b0000000001;
  assign MultLoop_acc_1205_nl = nl_MultLoop_acc_1205_nl[9:0];
  assign nl_MultLoop_acc_647_nl = (~ (data_rsci_idat[89:72])) + conv_s2s_17_18({(MultLoop_acc_1205_nl)
      , (data_rsci_idat[80:74])});
  assign MultLoop_acc_647_nl = nl_MultLoop_acc_647_nl[17:0];
  assign nl_MultLoop_acc_648_nl = ({(data_rsci_idat[89:72]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_647_nl);
  assign MultLoop_acc_648_nl = nl_MultLoop_acc_648_nl[19:0];
  assign nl_MultLoop_acc_649_nl = conv_s2s_23_24({(data_rsci_idat[89:72]) , 5'b00000})
      + conv_s2s_20_24(MultLoop_acc_648_nl);
  assign MultLoop_acc_649_nl = nl_MultLoop_acc_649_nl[23:0];
  assign nl_MultLoop_acc_1206_nl = conv_s2u_17_18(readslicef_24_17_7((MultLoop_acc_649_nl)))
      + (~ (data_rsci_idat[89:72]));
  assign MultLoop_acc_1206_nl = nl_MultLoop_acc_1206_nl[17:0];
  assign nl_MultLoop_acc_651_nl = conv_s2s_20_21({(data_rsci_idat[125:108]) , 2'b00})
      + conv_s2s_19_21(MultLoop_acc_650_cse_1);
  assign MultLoop_acc_651_nl = nl_MultLoop_acc_651_nl[20:0];
  assign nl_MultLoop_acc_349_nl = conv_s2u_21_24(MultLoop_acc_651_nl) + conv_s2u_23_24({(data_rsci_idat[125:108])
      , 5'b00000});
  assign MultLoop_acc_349_nl = nl_MultLoop_acc_349_nl[23:0];
  assign nl_MultLoop_acc_659_nl = (MultLoop_acc_657_nl) + (MultLoop_acc_1206_nl)
      + (readslicef_24_18_6((MultLoop_acc_349_nl)));
  assign MultLoop_acc_659_nl = nl_MultLoop_acc_659_nl[17:0];
  assign nl_MultLoop_acc_639_nl = ({(data_rsci_idat[107:90]) , 3'b001}) + conv_s2s_19_21({Result_Result_conc_60_18_7
      , (~ (data_rsci_idat[96:90]))});
  assign MultLoop_acc_639_nl = nl_MultLoop_acc_639_nl[20:0];
  assign nl_MultLoop_acc_640_nl = ({(~ (data_rsci_idat[107:90])) , 5'b00000}) + conv_s2s_21_23(MultLoop_acc_639_nl);
  assign MultLoop_acc_640_nl = nl_MultLoop_acc_640_nl[22:0];
  assign nl_MultLoop_acc_211_nl = conv_s2s_23_26(MultLoop_acc_640_nl) + conv_s2s_25_26({(~
      (data_rsci_idat[107:90])) , 7'b0100000});
  assign MultLoop_acc_211_nl = nl_MultLoop_acc_211_nl[25:0];
  assign nl_MultLoop_acc_205_nl = (MultLoop_acc_206_itm_20_4[16:1]) + 16'b0000000010001111;
  assign MultLoop_acc_205_nl = nl_MultLoop_acc_205_nl[15:0];
  assign nl_MultLoop_acc_635_nl = ({(data_rsci_idat[179:162]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_634_cse_1);
  assign MultLoop_acc_635_nl = nl_MultLoop_acc_635_nl[19:0];
  assign nl_MultLoop_acc_215_nl = conv_s2u_20_22(MultLoop_acc_635_nl) + ({(~ (data_rsci_idat[179:162]))
      , 4'b0000});
  assign MultLoop_acc_215_nl = nl_MultLoop_acc_215_nl[21:0];
  assign nl_MultLoop_acc_1207_nl = conv_s2s_11_12(data_rsci_idat[35:25]) + 12'b000000000001;
  assign MultLoop_acc_1207_nl = nl_MultLoop_acc_1207_nl[11:0];
  assign nl_MultLoop_acc_637_nl = conv_s2s_18_19(data_rsci_idat[35:18]) + conv_s2s_17_19({(MultLoop_acc_1207_nl)
      , (data_rsci_idat[24:20])});
  assign MultLoop_acc_637_nl = nl_MultLoop_acc_637_nl[18:0];
  assign nl_MultLoop_acc_207_nl = conv_s2u_19_23(MultLoop_acc_637_nl) + ({(~ (data_rsci_idat[35:18]))
      , 5'b00000});
  assign MultLoop_acc_207_nl = nl_MultLoop_acc_207_nl[22:0];
  assign nl_MultLoop_acc_632_nl = ({(data_rsci_idat[161:144]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[161:144]));
  assign MultLoop_acc_632_nl = nl_MultLoop_acc_632_nl[20:0];
  assign nl_MultLoop_acc_214_nl = conv_s2s_21_25(MultLoop_acc_632_nl) + conv_s2s_24_25({(data_rsci_idat[161:144])
      , 6'b000000});
  assign MultLoop_acc_214_nl = nl_MultLoop_acc_214_nl[24:0];
  assign nl_MultLoop_acc_658_nl = conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_211_nl)))
      + conv_s2s_17_18({(MultLoop_acc_205_nl) , (MultLoop_acc_206_itm_20_4[0])})
      + conv_s2s_15_18(readslicef_22_15_7((MultLoop_acc_215_nl))) + conv_s2s_15_18(MultLoop_acc_213_itm_22_7[15:1])
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_207_nl))) + conv_s2s_15_18(readslicef_25_15_10((MultLoop_acc_214_nl)));
  assign MultLoop_acc_658_nl = nl_MultLoop_acc_658_nl[17:0];
  assign nl_res_rsci_d_341_324  = (MultLoop_acc_659_nl) + (MultLoop_acc_658_nl);
  assign nl_MultLoop_acc_1199_nl = conv_s2u_16_17(MultLoop_acc_1198_itm_18_2[16:1])
      + (~ (data_rsci_idat[160:144]));
  assign MultLoop_acc_1199_nl = nl_MultLoop_acc_1199_nl[16:0];
  assign nl_MultLoop_acc_1201_nl = (~ (data_rsci_idat[179:162])) + conv_s2s_14_18(MultLoop_acc_777_sdt_1[19:6]);
  assign MultLoop_acc_1201_nl = nl_MultLoop_acc_1201_nl[17:0];
  assign nl_MultLoop_acc_1202_nl = conv_s2u_18_20(MultLoop_acc_1201_nl) + ({(data_rsci_idat[179:162])
      , 2'b01});
  assign MultLoop_acc_1202_nl = nl_MultLoop_acc_1202_nl[19:0];
  assign nl_MultLoop_acc_1200_nl =  -conv_s2s_14_15(data_rsci_idat[125:112]);
  assign MultLoop_acc_1200_nl = nl_MultLoop_acc_1200_nl[14:0];
  assign nl_MultLoop_acc_158_nl = conv_s2s_22_23({(~ (data_rsci_idat[125:108])) ,
      4'b0100}) + conv_s2s_20_23({(~ (data_rsci_idat[125:108])) , 2'b01}) + conv_s2s_19_23({(MultLoop_acc_1200_nl)
      , (~ (data_rsci_idat[111:108]))});
  assign MultLoop_acc_158_nl = nl_MultLoop_acc_158_nl[22:0];
  assign nl_MultLoop_acc_798_nl = conv_s2s_16_17(readslicef_20_16_4((MultLoop_acc_1202_nl)))
      + conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_158_nl))) + conv_s2s_15_17(MultLoop_acc_159_itm_24_9[15:1]);
  assign MultLoop_acc_798_nl = nl_MultLoop_acc_798_nl[16:0];
  assign nl_MultLoop_acc_801_nl = ({(MultLoop_acc_1199_nl) , (MultLoop_acc_1198_itm_18_2[0])})
      + conv_s2s_17_18(MultLoop_acc_798_nl);
  assign MultLoop_acc_801_nl = nl_MultLoop_acc_801_nl[17:0];
  assign nl_MultLoop_acc_1387_nl = conv_s2u_18_19(data_rsci_idat[107:90]) + conv_s2u_15_19(MultLoop_acc_753_cse_1[18:4]);
  assign MultLoop_acc_1387_nl = nl_MultLoop_acc_1387_nl[18:0];
  assign nl_MultLoop_acc_1192_nl = conv_s2u_17_18(readslicef_19_17_2((MultLoop_acc_1387_nl)))
      + (~ (data_rsci_idat[107:90]));
  assign MultLoop_acc_1192_nl = nl_MultLoop_acc_1192_nl[17:0];
  assign nl_MultLoop_acc_155_nl = conv_s2s_25_26({(~ (data_rsci_idat[71:54])) , 7'b0010000})
      + conv_s2s_22_26({(~ (data_rsci_idat[71:54])) , 4'b0001}) + conv_s2s_19_26({MultLoop_MultLoop_conc_202_18_7
      , (~ (data_rsci_idat[60:54]))});
  assign MultLoop_acc_155_nl = nl_MultLoop_acc_155_nl[25:0];
  assign nl_MultLoop_acc_1358_nl = conv_s2u_18_19(data_rsci_idat[89:72]) + conv_s2u_16_19(MultLoop_acc_786_cse_1[19:4]);
  assign MultLoop_acc_1358_nl = nl_MultLoop_acc_1358_nl[18:0];
  assign nl_MultLoop_acc_1194_nl = conv_s2u_16_19(readslicef_19_16_3((MultLoop_acc_1358_nl)))
      + conv_s2u_18_19(data_rsci_idat[89:72]);
  assign MultLoop_acc_1194_nl = nl_MultLoop_acc_1194_nl[18:0];
  assign nl_MultLoop_acc_790_nl = ({(data_rsci_idat[53:36]) , 4'b0100}) + conv_s2s_21_22(MultLoop_acc_789_cse_1);
  assign MultLoop_acc_790_nl = nl_MultLoop_acc_790_nl[21:0];
  assign nl_MultLoop_acc_791_nl = conv_s2s_24_25({(data_rsci_idat[53:36]) , 6'b000000})
      + conv_s2s_22_25(MultLoop_acc_790_nl);
  assign MultLoop_acc_791_nl = nl_MultLoop_acc_791_nl[24:0];
  assign nl_MultLoop_acc_1196_nl = conv_s2u_17_18(readslicef_25_17_8((MultLoop_acc_791_nl)))
      + (~ (data_rsci_idat[53:36]));
  assign MultLoop_acc_1196_nl = nl_MultLoop_acc_1196_nl[17:0];
  assign nl_MultLoop_acc_152_nl = conv_s2u_18_20(MultLoop_acc_412_cse_1) + ({(data_rsci_idat[17:0])
      , 2'b01});
  assign MultLoop_acc_152_nl = nl_MultLoop_acc_152_nl[19:0];
  assign nl_MultLoop_131_MultLoop_acc_3_nl = (readslicef_20_16_4((MultLoop_acc_152_nl)))
      + 16'b0000001100011001;
  assign MultLoop_131_MultLoop_acc_3_nl = nl_MultLoop_131_MultLoop_acc_3_nl[15:0];
  assign nl_MultLoop_acc_785_nl = (~ (data_rsci_idat[35:18])) + conv_s2s_13_18(data_rsci_idat[35:23]);
  assign MultLoop_acc_785_nl = nl_MultLoop_acc_785_nl[17:0];
  assign nl_MultLoop_acc_335_nl = conv_s2u_18_20(MultLoop_acc_785_nl) + ({(data_rsci_idat[35:18])
      , 2'b01});
  assign MultLoop_acc_335_nl = nl_MultLoop_acc_335_nl[19:0];
  assign nl_res_rsci_d_251_234  = (MultLoop_acc_801_nl) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_1192_nl)))
      + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_155_nl))) + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_1194_nl)))
      + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_1196_nl))) + conv_s2s_16_18(MultLoop_131_MultLoop_acc_3_nl)
      + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_335_nl)));
  assign nl_MultLoop_acc_669_nl = ({(data_rsci_idat[107:90]) , 4'b0001}) + conv_s2s_18_22(~
      (data_rsci_idat[107:90]));
  assign MultLoop_acc_669_nl = nl_MultLoop_acc_669_nl[21:0];
  assign nl_MultLoop_acc_1181_nl = conv_s2u_13_19(readslicef_22_13_9((MultLoop_acc_669_nl)))
      + conv_s2u_18_19(data_rsci_idat[107:90]);
  assign MultLoop_acc_1181_nl = nl_MultLoop_acc_1181_nl[18:0];
  assign nl_MultLoop_acc_1182_nl = conv_s2s_8_9(data_rsci_idat[125:118]) + 9'b000000001;
  assign MultLoop_acc_1182_nl = nl_MultLoop_acc_1182_nl[8:0];
  assign nl_MultLoop_acc_671_nl = (~ (data_rsci_idat[125:108])) + conv_s2s_17_18({(MultLoop_acc_1182_nl)
      , (data_rsci_idat[117:110])});
  assign MultLoop_acc_671_nl = nl_MultLoop_acc_671_nl[17:0];
  assign nl_MultLoop_acc_673_nl = ({(data_rsci_idat[125:108]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[125:108])) , 2'b01}) + conv_s2s_18_22(MultLoop_acc_671_nl);
  assign MultLoop_acc_673_nl = nl_MultLoop_acc_673_nl[21:0];
  assign nl_MultLoop_acc_674_nl = conv_s2s_24_25({(data_rsci_idat[125:108]) , 6'b000000})
      + conv_s2s_22_25(MultLoop_acc_673_nl);
  assign MultLoop_acc_674_nl = nl_MultLoop_acc_674_nl[24:0];
  assign nl_MultLoop_acc_1183_nl = conv_s2u_17_18(readslicef_25_17_8((MultLoop_acc_674_nl)))
      + (~ (data_rsci_idat[125:108]));
  assign MultLoop_acc_1183_nl = nl_MultLoop_acc_1183_nl[17:0];
  assign nl_MultLoop_acc_677_nl = conv_s2s_26_27({(~ (data_rsci_idat[161:144])) ,
      8'b01000000}) + conv_s2s_24_27({(~ (data_rsci_idat[161:144])) , 6'b010000})
      + conv_s2s_22_27({(~ (data_rsci_idat[161:144])) , 4'b0001}) + conv_s2s_18_27(~
      (data_rsci_idat[161:144]));
  assign MultLoop_acc_677_nl = nl_MultLoop_acc_677_nl[26:0];
  assign nl_MultLoop_acc_1184_nl = conv_s2u_19_20(readslicef_27_19_8((MultLoop_acc_677_nl)))
      + ({(data_rsci_idat[161:144]) , 2'b01});
  assign MultLoop_acc_1184_nl = nl_MultLoop_acc_1184_nl[19:0];
  assign nl_MultLoop_acc_1356_nl = conv_s2u_18_19(data_rsci_idat[179:162]) + conv_s2u_16_19(MultLoop_acc_702_cse_1[18:3]);
  assign MultLoop_acc_1356_nl = nl_MultLoop_acc_1356_nl[18:0];
  assign nl_MultLoop_acc_1185_nl = conv_s2u_15_19(readslicef_19_15_4((MultLoop_acc_1356_nl)))
      + conv_s2u_18_19(data_rsci_idat[179:162]);
  assign MultLoop_acc_1185_nl = nl_MultLoop_acc_1185_nl[18:0];
  assign nl_MultLoop_acc_687_nl = (readslicef_19_18_1((MultLoop_acc_1181_nl))) +
      (MultLoop_acc_1183_nl) + (readslicef_20_18_2((MultLoop_acc_1184_nl))) + (readslicef_19_18_1((MultLoop_acc_1185_nl)));
  assign MultLoop_acc_687_nl = nl_MultLoop_acc_687_nl[17:0];
  assign nl_MultLoop_acc_663_nl = ({(data_rsci_idat[35:18]) , 4'b0001}) + conv_s2s_19_22({MultLoop_MultLoop_conc_210_18_8
      , (~ (data_rsci_idat[25:18]))});
  assign MultLoop_acc_663_nl = nl_MultLoop_acc_663_nl[21:0];
  assign nl_MultLoop_acc_664_nl = conv_s2s_24_25({(data_rsci_idat[35:18]) , 6'b000000})
      + conv_s2s_22_25(MultLoop_acc_663_nl);
  assign MultLoop_acc_664_nl = nl_MultLoop_acc_664_nl[24:0];
  assign nl_MultLoop_acc_1187_nl = conv_s2u_17_18(readslicef_25_17_8((MultLoop_acc_664_nl)))
      + (~ (data_rsci_idat[35:18]));
  assign MultLoop_acc_1187_nl = nl_MultLoop_acc_1187_nl[17:0];
  assign nl_MultLoop_acc_194_nl = conv_s2u_15_18(data_rsci_idat[17:3]) - (data_rsci_idat[17:0]);
  assign MultLoop_acc_194_nl = nl_MultLoop_acc_194_nl[17:0];
  assign nl_MultLoop_171_MultLoop_acc_3_nl = (readslicef_18_15_3((MultLoop_acc_194_nl)))
      + 15'b111110111110111;
  assign MultLoop_171_MultLoop_acc_3_nl = nl_MultLoop_171_MultLoop_acc_3_nl[14:0];
  assign nl_MultLoop_acc_680_nl = conv_s2s_15_16(MultLoop_171_MultLoop_acc_3_nl)
      + conv_s2s_12_16(Result_acc_175_cse[18:7]);
  assign MultLoop_acc_680_nl = nl_MultLoop_acc_680_nl[15:0];
  assign nl_MultLoop_acc_682_nl = (readslicef_18_17_1((MultLoop_acc_1187_nl))) +
      conv_s2s_16_17(MultLoop_acc_680_nl);
  assign MultLoop_acc_682_nl = nl_MultLoop_acc_682_nl[16:0];
  assign nl_MultLoop_acc_1357_nl = conv_s2u_19_22(MultLoop_acc_660_itm_22_4_1) +
      ({(data_rsci_idat[89:72]) , 4'b0001});
  assign MultLoop_acc_1357_nl = nl_MultLoop_acc_1357_nl[21:0];
  assign nl_MultLoop_acc_661_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_13_18(data_rsci_idat[53:41]);
  assign MultLoop_acc_661_nl = nl_MultLoop_acc_661_nl[17:0];
  assign nl_MultLoop_acc_346_nl = conv_s2u_18_21(MultLoop_acc_661_nl) + ({(data_rsci_idat[53:36])
      , 3'b001});
  assign MultLoop_acc_346_nl = nl_MultLoop_acc_346_nl[20:0];
  assign nl_MultLoop_acc_683_nl = conv_s2s_17_18(MultLoop_acc_682_nl) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1357_nl)))
      + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_346_nl)));
  assign MultLoop_acc_683_nl = nl_MultLoop_acc_683_nl[17:0];
  assign nl_MultLoop_acc_667_nl = ({(data_rsci_idat[71:54]) , 5'b01000}) + conv_s2s_21_23({(~
      (data_rsci_idat[71:54])) , 3'b001}) + conv_s2s_19_23({MultLoop_MultLoop_conc_228_18_9
      , (~ (data_rsci_idat[62:54]))});
  assign MultLoop_acc_667_nl = nl_MultLoop_acc_667_nl[22:0];
  assign nl_MultLoop_acc_1189_nl = (~ (data_rsci_idat[71:54])) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_667_nl)));
  assign MultLoop_acc_1189_nl = nl_MultLoop_acc_1189_nl[17:0];
  assign nl_MultLoop_acc_1190_nl = conv_s2u_18_21(MultLoop_acc_1189_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[71:54])) , 2'b01});
  assign MultLoop_acc_1190_nl = nl_MultLoop_acc_1190_nl[20:0];
  assign nl_MultLoop_acc_686_nl = (MultLoop_acc_683_nl) + (readslicef_21_18_3((MultLoop_acc_1190_nl)));
  assign MultLoop_acc_686_nl = nl_MultLoop_acc_686_nl[17:0];
  assign nl_res_rsci_d_323_306  = (MultLoop_acc_687_nl) + (MultLoop_acc_686_nl);
  assign nl_MultLoop_acc_1172_nl = (~ (data_rsci_idat[35:18])) + conv_s2s_15_18(MultLoop_acc_759_sdt_1[20:6]);
  assign MultLoop_acc_1172_nl = nl_MultLoop_acc_1172_nl[17:0];
  assign nl_MultLoop_acc_1352_nl = conv_s2u_20_21({(~ (data_rsci_idat[35:18])) ,
      2'b01}) + conv_s2u_18_21(MultLoop_acc_1172_nl);
  assign MultLoop_acc_1352_nl = nl_MultLoop_acc_1352_nl[20:0];
  assign nl_MultLoop_acc_1173_nl = conv_s2u_19_20(readslicef_21_19_2((MultLoop_acc_1352_nl)))
      + ({(data_rsci_idat[35:18]) , 2'b01});
  assign MultLoop_acc_1173_nl = nl_MultLoop_acc_1173_nl[19:0];
  assign nl_MultLoop_acc_764_nl = ({(data_rsci_idat[161:144]) , 4'b0100}) + conv_s2s_21_22(MultLoop_acc_763_cse_1);
  assign MultLoop_acc_764_nl = nl_MultLoop_acc_764_nl[21:0];
  assign nl_MultLoop_acc_765_nl = conv_s2s_24_25({(data_rsci_idat[161:144]) , 6'b000000})
      + conv_s2s_22_25(MultLoop_acc_764_nl);
  assign MultLoop_acc_765_nl = nl_MultLoop_acc_765_nl[24:0];
  assign nl_MultLoop_acc_1175_nl = conv_s2u_17_18(readslicef_25_17_8((MultLoop_acc_765_nl)))
      + (~ (data_rsci_idat[161:144]));
  assign MultLoop_acc_1175_nl = nl_MultLoop_acc_1175_nl[17:0];
  assign nl_MultLoop_acc_772_nl = (readslicef_20_18_2((MultLoop_acc_1173_nl))) +
      (MultLoop_acc_1175_nl);
  assign MultLoop_acc_772_nl = nl_MultLoop_acc_772_nl[17:0];
  assign nl_MultLoop_acc_749_nl = ({(~ (data_rsci_idat[179:162])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[179:162])
      + conv_s2s_17_20({MultLoop_MultLoop_conc_224_16_6 , (data_rsci_idat[169:164])});
  assign MultLoop_acc_749_nl = nl_MultLoop_acc_749_nl[19:0];
  assign nl_MultLoop_acc_750_nl = conv_s2s_22_23({(~ (data_rsci_idat[179:162])) ,
      4'b0100}) + conv_s2s_20_23(MultLoop_acc_749_nl);
  assign MultLoop_acc_750_nl = nl_MultLoop_acc_750_nl[22:0];
  assign nl_MultLoop_acc_339_nl = conv_s2u_23_25(MultLoop_acc_750_nl) + conv_s2u_24_25({(~
      (data_rsci_idat[179:162])) , 6'b010000});
  assign MultLoop_acc_339_nl = nl_MultLoop_acc_339_nl[24:0];
  assign nl_MultLoop_acc_1353_nl = conv_s2u_16_19(MultLoop_acc_751_itm_18_2[16:1])
      + conv_s2u_18_19(data_rsci_idat[125:108]);
  assign MultLoop_acc_1353_nl = nl_MultLoop_acc_1353_nl[18:0];
  assign nl_MultLoop_acc_771_nl = conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_339_nl)))
      + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_1353_nl)));
  assign MultLoop_acc_771_nl = nl_MultLoop_acc_771_nl[17:0];
  assign nl_MultLoop_acc_774_nl = (MultLoop_acc_772_nl) + (MultLoop_acc_771_nl);
  assign MultLoop_acc_774_nl = nl_MultLoop_acc_774_nl[17:0];
  assign nl_MultLoop_acc_754_nl = ({(~ (data_rsci_idat[107:90])) , 4'b0000}) + conv_s2s_19_22(MultLoop_acc_753_cse_1);
  assign MultLoop_acc_754_nl = nl_MultLoop_acc_754_nl[21:0];
  assign nl_MultLoop_acc_337_nl = conv_s2u_22_25(MultLoop_acc_754_nl) + conv_s2u_24_25({(~
      (data_rsci_idat[107:90])) , 6'b010000});
  assign MultLoop_acc_337_nl = nl_MultLoop_acc_337_nl[24:0];
  assign nl_MultLoop_acc_756_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_17_18({MultLoop_acc_1178_cse_1
      , (data_rsci_idat[41:38])});
  assign MultLoop_acc_756_nl = nl_MultLoop_acc_756_nl[17:0];
  assign nl_MultLoop_acc_757_nl = ({(data_rsci_idat[53:36]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_756_nl);
  assign MultLoop_acc_757_nl = nl_MultLoop_acc_757_nl[19:0];
  assign nl_MultLoop_acc_165_nl = conv_s2u_20_22(MultLoop_acc_757_nl) + ({(~ (data_rsci_idat[53:36]))
      , 4'b0000});
  assign MultLoop_acc_165_nl = nl_MultLoop_acc_165_nl[21:0];
  assign nl_MultLoop_acc_758_nl = (~ (data_rsci_idat[71:54])) + conv_s2s_11_18(data_rsci_idat[71:61]);
  assign MultLoop_acc_758_nl = nl_MultLoop_acc_758_nl[17:0];
  assign nl_MultLoop_acc_336_nl = conv_s2u_18_20(MultLoop_acc_758_nl) + ({(data_rsci_idat[71:54])
      , 2'b01});
  assign MultLoop_acc_336_nl = nl_MultLoop_acc_336_nl[19:0];
  assign nl_MultLoop_acc_1179_nl = conv_s2u_15_19(MultLoop_acc_1354_itm_19_3[16:2])
      + conv_s2u_18_19(data_rsci_idat[89:72]);
  assign MultLoop_acc_1179_nl = nl_MultLoop_acc_1179_nl[18:0];
  assign nl_MultLoop_acc_1355_nl = conv_s2u_19_21(MultLoop_acc_744_cse_1[20:2]) +
      ({(data_rsci_idat[17:0]) , 3'b001});
  assign MultLoop_acc_1355_nl = nl_MultLoop_acc_1355_nl[20:0];
  assign nl_MultLoop_acc_1180_nl = conv_s2u_8_9(MultLoop_acc_170_itm_17_8[9:2]) +
      9'b011111011;
  assign MultLoop_acc_1180_nl = nl_MultLoop_acc_1180_nl[8:0];
  assign nl_MultLoop_acc_767_nl = conv_s2s_13_14(readslicef_21_13_8((MultLoop_acc_1355_nl)))
      + conv_u2s_11_14({(MultLoop_acc_1180_nl) , (MultLoop_acc_170_itm_17_8[1:0])});
  assign MultLoop_acc_767_nl = nl_MultLoop_acc_767_nl[13:0];
  assign nl_MultLoop_acc_768_nl = (readslicef_19_16_3((MultLoop_acc_1179_nl))) +
      conv_s2s_14_16(MultLoop_acc_767_nl);
  assign MultLoop_acc_768_nl = nl_MultLoop_acc_768_nl[15:0];
  assign nl_res_rsci_d_269_252  = (MultLoop_acc_774_nl) + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_337_nl)))
      + conv_s2s_17_18(readslicef_22_17_5((MultLoop_acc_165_nl))) + conv_s2s_17_18(readslicef_20_17_3((MultLoop_acc_336_nl)))
      + conv_s2s_16_18(MultLoop_acc_768_nl);
  assign nl_MultLoop_acc_696_nl = ({(data_rsci_idat[53:36]) , 7'b0100000}) + conv_s2s_23_25({(~
      (data_rsci_idat[53:36])) , 5'b00001}) + conv_s2s_18_25(~ (data_rsci_idat[53:36]));
  assign MultLoop_acc_696_nl = nl_MultLoop_acc_696_nl[24:0];
  assign nl_MultLoop_acc_1165_nl = conv_s2u_16_19(readslicef_25_16_9((MultLoop_acc_696_nl)))
      + conv_s2u_18_19(data_rsci_idat[53:36]);
  assign MultLoop_acc_1165_nl = nl_MultLoop_acc_1165_nl[18:0];
  assign nl_MultLoop_acc_697_nl = (~ (data_rsci_idat[107:90])) + conv_s2s_16_18(data_rsci_idat[107:92]);
  assign MultLoop_acc_697_nl = nl_MultLoop_acc_697_nl[17:0];
  assign nl_MultLoop_acc_698_nl = ({(data_rsci_idat[107:90]) , 4'b0001}) + conv_s2s_18_22(MultLoop_acc_697_nl);
  assign MultLoop_acc_698_nl = nl_MultLoop_acc_698_nl[21:0];
  assign nl_MultLoop_acc_1166_nl = conv_s2u_15_19(readslicef_22_15_7((MultLoop_acc_698_nl)))
      + conv_s2u_18_19(data_rsci_idat[107:90]);
  assign MultLoop_acc_1166_nl = nl_MultLoop_acc_1166_nl[18:0];
  assign nl_MultLoop_acc_1167_nl = conv_s2s_10_11(data_rsci_idat[125:116]) + 11'b00000000001;
  assign MultLoop_acc_1167_nl = nl_MultLoop_acc_1167_nl[10:0];
  assign nl_MultLoop_acc_701_nl = ({(~ (data_rsci_idat[125:108])) , 3'b000}) + conv_s2s_18_21(data_rsci_idat[125:108])
      + conv_s2s_16_21({(MultLoop_acc_1167_nl) , (data_rsci_idat[115:111])});
  assign MultLoop_acc_701_nl = nl_MultLoop_acc_701_nl[20:0];
  assign nl_MultLoop_acc_343_nl = conv_s2u_21_24(MultLoop_acc_701_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[125:108])) , 5'b01000});
  assign MultLoop_acc_343_nl = nl_MultLoop_acc_343_nl[23:0];
  assign nl_MultLoop_acc_1168_nl = conv_s2u_14_19(MultLoop_acc_1350_itm_18_5) + conv_s2u_18_19(data_rsci_idat[179:162]);
  assign MultLoop_acc_1168_nl = nl_MultLoop_acc_1168_nl[18:0];
  assign nl_MultLoop_acc_712_nl = (readslicef_19_18_1((MultLoop_acc_1165_nl))) +
      (readslicef_19_18_1((MultLoop_acc_1166_nl))) + (readslicef_24_18_6((MultLoop_acc_343_nl)))
      + (readslicef_19_18_1((MultLoop_acc_1168_nl)));
  assign MultLoop_acc_712_nl = nl_MultLoop_acc_712_nl[17:0];
  assign nl_MultLoop_acc_1169_nl = conv_s2s_11_12(data_rsci_idat[143:133]) + 12'b000000000001;
  assign MultLoop_acc_1169_nl = nl_MultLoop_acc_1169_nl[11:0];
  assign nl_MultLoop_acc_691_nl = (~ (data_rsci_idat[143:126])) + conv_s2s_14_18({(MultLoop_acc_1169_nl)
      , (data_rsci_idat[132:131])});
  assign MultLoop_acc_691_nl = nl_MultLoop_acc_691_nl[17:0];
  assign nl_MultLoop_acc_344_nl = conv_s2u_18_21(MultLoop_acc_691_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[143:126])) , 2'b01});
  assign MultLoop_acc_344_nl = nl_MultLoop_acc_344_nl[20:0];
  assign nl_MultLoop_acc_188_nl = conv_s2s_19_25({Result_Result_conc_56_18_6 , (~
      (data_rsci_idat[77:72]))}) + conv_s2s_24_25({(~ (data_rsci_idat[89:72])) ,
      6'b000001});
  assign MultLoop_acc_188_nl = nl_MultLoop_acc_188_nl[24:0];
  assign nl_MultLoop_acc_1351_nl = conv_s2u_18_21(MultLoop_acc_694_itm_19_2_1) +
      ({(data_rsci_idat[71:54]) , 3'b001});
  assign MultLoop_acc_1351_nl = nl_MultLoop_acc_1351_nl[20:0];
  assign nl_MultLoop_acc_185_nl = conv_s2u_12_18(data_rsci_idat[35:24]) - (data_rsci_idat[35:18]);
  assign MultLoop_acc_185_nl = nl_MultLoop_acc_185_nl[17:0];
  assign nl_MultLoop_acc_704_nl = conv_s2s_14_15(readslicef_18_14_4((MultLoop_acc_185_nl)))
      + 15'b000000010001011;
  assign MultLoop_acc_704_nl = nl_MultLoop_acc_704_nl[14:0];
  assign nl_MultLoop_acc_184_nl = conv_s2s_23_24({(~ (data_rsci_idat[17:0])) , 5'b01000})
      + conv_s2s_21_24({(~ (data_rsci_idat[17:0])) , 3'b001}) + conv_s2s_19_24({MultLoop_MultLoop_conc_206_18_5
      , (~ (data_rsci_idat[4:0]))});
  assign MultLoop_acc_184_nl = nl_MultLoop_acc_184_nl[23:0];
  assign nl_MultLoop_acc_711_nl = conv_s2s_17_18(readslicef_21_17_4((MultLoop_acc_344_nl)))
      + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_188_nl))) + conv_s2s_17_18(readslicef_21_17_4((MultLoop_acc_1351_nl)))
      + conv_s2s_15_18(MultLoop_acc_704_nl) + conv_s2s_14_18(MultLoop_acc_108_itm_19_6)
      + conv_s2s_14_18(readslicef_24_14_10((MultLoop_acc_184_nl)));
  assign MultLoop_acc_711_nl = nl_MultLoop_acc_711_nl[17:0];
  assign nl_res_rsci_d_305_288  = (MultLoop_acc_712_nl) + (MultLoop_acc_711_nl);
  assign nl_MultLoop_acc_179_nl = conv_s2s_24_25({(~ (data_rsci_idat[107:90])) ,
      6'b001000}) + conv_s2s_21_25({(~ (data_rsci_idat[107:90])) , 3'b001}) + conv_s2s_19_25({Result_Result_conc_62_18_6
      , (~ (data_rsci_idat[95:90]))});
  assign MultLoop_acc_179_nl = nl_MultLoop_acc_179_nl[24:0];
  assign nl_MultLoop_acc_1162_nl =  -conv_s2s_12_13(data_rsci_idat[35:24]);
  assign MultLoop_acc_1162_nl = nl_MultLoop_acc_1162_nl[12:0];
  assign nl_MultLoop_acc_730_nl = ({(data_rsci_idat[35:18]) , 4'b0001}) + conv_s2s_19_22({(MultLoop_acc_1162_nl)
      , (~ (data_rsci_idat[23:18]))});
  assign MultLoop_acc_730_nl = nl_MultLoop_acc_730_nl[21:0];
  assign nl_MultLoop_acc_1163_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_730_nl)))
      + (~ (data_rsci_idat[35:18]));
  assign MultLoop_acc_1163_nl = nl_MultLoop_acc_1163_nl[17:0];
  assign nl_MultLoop_acc_732_nl = (readslicef_18_14_4((MultLoop_acc_1163_nl))) +
      14'b11111111011101;
  assign MultLoop_acc_732_nl = nl_MultLoop_acc_732_nl[13:0];
  assign nl_MultLoop_acc_1349_nl = conv_s2u_14_19(MultLoop_acc_731_itm_18_4[14:1])
      + conv_s2u_18_19(data_rsci_idat[17:0]);
  assign MultLoop_acc_1349_nl = nl_MultLoop_acc_1349_nl[18:0];
  assign nl_MultLoop_152_MultLoop_acc_3_nl = conv_s2s_14_17(MultLoop_acc_732_nl)
      + (readslicef_19_17_2((MultLoop_acc_1349_nl)));
  assign MultLoop_152_MultLoop_acc_3_nl = nl_MultLoop_152_MultLoop_acc_3_nl[16:0];
  assign nl_MultLoop_acc_734_nl = ({(~ (data_rsci_idat[53:36])) , 4'b0000}) + conv_s2s_20_22(MultLoop_acc_733_cse_1);
  assign MultLoop_acc_734_nl = nl_MultLoop_acc_734_nl[21:0];
  assign nl_MultLoop_acc_735_nl = ({(data_rsci_idat[53:36]) , 6'b010000}) + conv_s2s_22_24(MultLoop_acc_734_nl);
  assign MultLoop_acc_735_nl = nl_MultLoop_acc_735_nl[23:0];
  assign nl_MultLoop_acc_1164_nl = conv_s2u_16_19(readslicef_24_16_8((MultLoop_acc_735_nl)))
      + conv_s2u_18_19(data_rsci_idat[53:36]);
  assign MultLoop_acc_1164_nl = nl_MultLoop_acc_1164_nl[18:0];
  assign nl_MultLoop_acc_340_nl = conv_s2u_18_23(MultLoop_acc_410_cse_1) + ({(data_rsci_idat[71:54])
      , 5'b00001});
  assign MultLoop_acc_340_nl = nl_MultLoop_acc_340_nl[22:0];
  assign nl_MultLoop_acc_742_nl = conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_179_nl)))
      + conv_s2s_17_18(MultLoop_152_MultLoop_acc_3_nl) + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_1164_nl)))
      + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_340_nl)));
  assign MultLoop_acc_742_nl = nl_MultLoop_acc_742_nl[17:0];
  assign nl_MultLoop_acc_718_nl = ({(data_rsci_idat[179:162]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[179:162])) , 2'b01}) + conv_s2s_19_22({MultLoop_MultLoop_conc_216_18_8
      , (~ (data_rsci_idat[169:162]))});
  assign MultLoop_acc_718_nl = nl_MultLoop_acc_718_nl[21:0];
  assign nl_MultLoop_acc_719_nl = conv_s2s_24_25({(data_rsci_idat[179:162]) , 6'b000000})
      + conv_s2s_22_25(MultLoop_acc_718_nl);
  assign MultLoop_acc_719_nl = nl_MultLoop_acc_719_nl[24:0];
  assign nl_MultLoop_acc_1155_nl = conv_s2u_17_18(readslicef_25_17_8((MultLoop_acc_719_nl)))
      + (~ (data_rsci_idat[179:162]));
  assign MultLoop_acc_1155_nl = nl_MultLoop_acc_1155_nl[17:0];
  assign nl_MultLoop_acc_1386_nl = conv_s2u_18_19(data_rsci_idat[161:144]) + conv_s2u_14_19(MultLoop_acc_714_itm_19_4[15:2]);
  assign MultLoop_acc_1386_nl = nl_MultLoop_acc_1386_nl[18:0];
  assign nl_MultLoop_acc_1153_nl = conv_s2u_17_18(readslicef_19_17_2((MultLoop_acc_1386_nl)))
      + (~ (data_rsci_idat[161:144]));
  assign MultLoop_acc_1153_nl = nl_MultLoop_acc_1153_nl[17:0];
  assign nl_MultLoop_acc_722_nl = ({(data_rsci_idat[125:108]) , 7'b0100000}) + conv_s2s_23_25({(~
      (data_rsci_idat[125:108])) , 5'b00001}) + conv_s2s_19_25({MultLoop_MultLoop_conc_222_18_9
      , (~ (data_rsci_idat[116:108]))});
  assign MultLoop_acc_722_nl = nl_MultLoop_acc_722_nl[24:0];
  assign nl_MultLoop_acc_1157_nl = conv_s2u_16_18(readslicef_25_16_9((MultLoop_acc_722_nl)))
      + (~ (data_rsci_idat[125:108]));
  assign MultLoop_acc_1157_nl = nl_MultLoop_acc_1157_nl[17:0];
  assign nl_MultLoop_acc_724_nl = ({(data_rsci_idat[89:72]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_204_18_9
      , (~ (data_rsci_idat[80:72]))});
  assign MultLoop_acc_724_nl = nl_MultLoop_acc_724_nl[19:0];
  assign nl_MultLoop_acc_725_nl = conv_s2s_22_23({(data_rsci_idat[89:72]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_724_nl);
  assign MultLoop_acc_725_nl = nl_MultLoop_acc_725_nl[22:0];
  assign nl_MultLoop_acc_1159_nl = conv_s2u_18_19(data_rsci_idat[89:72]) + conv_s2u_16_19(readslicef_23_16_7((MultLoop_acc_725_nl)));
  assign MultLoop_acc_1159_nl = nl_MultLoop_acc_1159_nl[18:0];
  assign nl_MultLoop_acc_1160_nl = conv_s2u_17_18(readslicef_19_17_2((MultLoop_acc_1159_nl)))
      + (~ (data_rsci_idat[89:72]));
  assign MultLoop_acc_1160_nl = nl_MultLoop_acc_1160_nl[17:0];
  assign nl_res_rsci_d_287_270  = (MultLoop_acc_742_nl) + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_1155_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_1153_nl))) + conv_s2s_16_18(MultLoop_acc_159_itm_24_9)
      + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_1157_nl))) + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_1160_nl)));

  function automatic [9:0] readslicef_18_10_8;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_18_10_8 = tmp[9:0];
  end
  endfunction


  function automatic [10:0] readslicef_18_11_7;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_18_11_7 = tmp[10:0];
  end
  endfunction


  function automatic [11:0] readslicef_18_12_6;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_18_12_6 = tmp[11:0];
  end
  endfunction


  function automatic [13:0] readslicef_18_14_4;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_18_14_4 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_18_15_3;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_18_15_3 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_18_16_2;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_18_16_2 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_18_17_1;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_18_17_1 = tmp[16:0];
  end
  endfunction


  function automatic [12:0] readslicef_19_13_6;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_19_13_6 = tmp[12:0];
  end
  endfunction


  function automatic [13:0] readslicef_19_14_5;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_19_14_5 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_19_15_4;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_19_15_4 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_19_16_3;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_19_16_3 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_19_17_2;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_19_17_2 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_19_18_1;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_19_18_1 = tmp[17:0];
  end
  endfunction


  function automatic [10:0] readslicef_20_11_9;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_20_11_9 = tmp[10:0];
  end
  endfunction


  function automatic [11:0] readslicef_20_12_8;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_20_12_8 = tmp[11:0];
  end
  endfunction


  function automatic [12:0] readslicef_20_13_7;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_20_13_7 = tmp[12:0];
  end
  endfunction


  function automatic [13:0] readslicef_20_14_6;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_20_14_6 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_20_15_5;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_20_15_5 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_20_16_4;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_20_16_4 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_20_17_3;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_20_17_3 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_20_18_2;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_20_18_2 = tmp[17:0];
  end
  endfunction


  function automatic [10:0] readslicef_21_11_10;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_21_11_10 = tmp[10:0];
  end
  endfunction


  function automatic [12:0] readslicef_21_13_8;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_21_13_8 = tmp[12:0];
  end
  endfunction


  function automatic [13:0] readslicef_21_14_7;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_21_14_7 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_21_15_6;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_21_15_6 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_21_16_5;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_21_16_5 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_21_17_4;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_21_17_4 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_21_18_3;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_21_18_3 = tmp[17:0];
  end
  endfunction


  function automatic [18:0] readslicef_21_19_2;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_21_19_2 = tmp[18:0];
  end
  endfunction


  function automatic [11:0] readslicef_22_12_10;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_22_12_10 = tmp[11:0];
  end
  endfunction


  function automatic [12:0] readslicef_22_13_9;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_22_13_9 = tmp[12:0];
  end
  endfunction


  function automatic [13:0] readslicef_22_14_8;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_22_14_8 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_22_15_7;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_22_15_7 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_22_16_6;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_22_16_6 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_22_17_5;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_22_17_5 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_22_18_4;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_22_18_4 = tmp[17:0];
  end
  endfunction


  function automatic [18:0] readslicef_22_19_3;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_22_19_3 = tmp[18:0];
  end
  endfunction


  function automatic [12:0] readslicef_23_13_10;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_23_13_10 = tmp[12:0];
  end
  endfunction


  function automatic [13:0] readslicef_23_14_9;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_23_14_9 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_23_15_8;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_23_15_8 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_23_16_7;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_23_16_7 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_23_17_6;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_23_17_6 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_23_18_5;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_23_18_5 = tmp[17:0];
  end
  endfunction


  function automatic [18:0] readslicef_23_19_4;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_23_19_4 = tmp[18:0];
  end
  endfunction


  function automatic [13:0] readslicef_24_14_10;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_24_14_10 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_24_15_9;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_24_15_9 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_24_16_8;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_24_16_8 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_24_17_7;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_24_17_7 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_24_18_6;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_24_18_6 = tmp[17:0];
  end
  endfunction


  function automatic [18:0] readslicef_24_19_5;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_24_19_5 = tmp[18:0];
  end
  endfunction


  function automatic [14:0] readslicef_25_15_10;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_25_15_10 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_25_16_9;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_25_16_9 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_25_17_8;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_25_17_8 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_25_18_7;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_25_18_7 = tmp[17:0];
  end
  endfunction


  function automatic [15:0] readslicef_26_16_10;
    input [25:0] vector;
    reg [25:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_26_16_10 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_26_17_9;
    input [25:0] vector;
    reg [25:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_26_17_9 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_26_18_8;
    input [25:0] vector;
    reg [25:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_26_18_8 = tmp[17:0];
  end
  endfunction


  function automatic [18:0] readslicef_26_19_7;
    input [25:0] vector;
    reg [25:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_26_19_7 = tmp[18:0];
  end
  endfunction


  function automatic [16:0] readslicef_27_17_10;
    input [26:0] vector;
    reg [26:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_27_17_10 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_27_18_9;
    input [26:0] vector;
    reg [26:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_27_18_9 = tmp[17:0];
  end
  endfunction


  function automatic [18:0] readslicef_27_19_8;
    input [26:0] vector;
    reg [26:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_27_19_8 = tmp[18:0];
  end
  endfunction


  function automatic [17:0] readslicef_28_18_10;
    input [27:0] vector;
    reg [27:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_28_18_10 = tmp[17:0];
  end
  endfunction


  function automatic [8:0] conv_s2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_9 = {vector[7], vector};
  end
  endfunction


  function automatic [9:0] conv_s2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_10 = {vector[8], vector};
  end
  endfunction


  function automatic [10:0] conv_s2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_s2s_10_11 = {vector[9], vector};
  end
  endfunction


  function automatic [11:0] conv_s2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_12 = {vector[10], vector};
  end
  endfunction


  function automatic [13:0] conv_s2s_11_14 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_14 = {{3{vector[10]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_11_18 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_18 = {{7{vector[10]}}, vector};
  end
  endfunction


  function automatic [12:0] conv_s2s_12_13 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_13 = {vector[11], vector};
  end
  endfunction


  function automatic [13:0] conv_s2s_12_14 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_14 = {{2{vector[11]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_12_16 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_16 = {{4{vector[11]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_12_17 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_17 = {{5{vector[11]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_12_18 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_18 = {{6{vector[11]}}, vector};
  end
  endfunction


  function automatic [13:0] conv_s2s_13_14 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_14 = {vector[12], vector};
  end
  endfunction


  function automatic [14:0] conv_s2s_13_15 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_15 = {{2{vector[12]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_13_17 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_17 = {{4{vector[12]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_13_18 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_18 = {{5{vector[12]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_13_19 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_19 = {{6{vector[12]}}, vector};
  end
  endfunction


  function automatic [14:0] conv_s2s_14_15 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_15 = {vector[13], vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_14_16 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_16 = {{2{vector[13]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_14_17 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_17 = {{3{vector[13]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_14_18 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_18 = {{4{vector[13]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_14_19 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_19 = {{5{vector[13]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_15_16 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_16 = {vector[14], vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_15_17 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_17 = {{2{vector[14]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_15_18 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_18 = {{3{vector[14]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_15_19 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_19 = {{4{vector[14]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_15_20 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_20 = {{5{vector[14]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_15_21 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_21 = {{6{vector[14]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_16_17 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_17 = {vector[15], vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_16_18 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_18 = {{2{vector[15]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_16_19 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_19 = {{3{vector[15]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_16_20 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_20 = {{4{vector[15]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_16_21 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_21 = {{5{vector[15]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_17_18 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_18 = {vector[16], vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_17_19 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_19 = {{2{vector[16]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_17_20 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_20 = {{3{vector[16]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_17_21 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_21 = {{4{vector[16]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_17_22 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_22 = {{5{vector[16]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_17_23 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_23 = {{6{vector[16]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_19 = {vector[17], vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_18_20 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_20 = {{2{vector[17]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_18_21 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_21 = {{3{vector[17]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_18_22 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_22 = {{4{vector[17]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_18_23 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_23 = {{5{vector[17]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_18_24 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_24 = {{6{vector[17]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_18_25 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_25 = {{7{vector[17]}}, vector};
  end
  endfunction


  function automatic [26:0] conv_s2s_18_27 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_27 = {{9{vector[17]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_19_20 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_20 = {vector[18], vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_19_21 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_21 = {{2{vector[18]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_19_22 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_22 = {{3{vector[18]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_19_23 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_23 = {{4{vector[18]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_19_24 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_24 = {{5{vector[18]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_19_25 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_25 = {{6{vector[18]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_19_26 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_26 = {{7{vector[18]}}, vector};
  end
  endfunction


  function automatic [26:0] conv_s2s_19_27 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_27 = {{8{vector[18]}}, vector};
  end
  endfunction


  function automatic [27:0] conv_s2s_19_28 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_28 = {{9{vector[18]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_20_21 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_21 = {vector[19], vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_20_22 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_22 = {{2{vector[19]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_20_23 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_23 = {{3{vector[19]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_20_24 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_24 = {{4{vector[19]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_20_25 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_25 = {{5{vector[19]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_20_26 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_26 = {{6{vector[19]}}, vector};
  end
  endfunction


  function automatic [26:0] conv_s2s_20_27 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_27 = {{7{vector[19]}}, vector};
  end
  endfunction


  function automatic [27:0] conv_s2s_20_28 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_28 = {{8{vector[19]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_21_22 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_22 = {vector[20], vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_21_23 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_23 = {{2{vector[20]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_21_24 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_24 = {{3{vector[20]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_21_25 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_25 = {{4{vector[20]}}, vector};
  end
  endfunction


  function automatic [26:0] conv_s2s_21_27 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_27 = {{6{vector[20]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_22_23 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_23 = {vector[21], vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_22_24 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_24 = {{2{vector[21]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_22_25 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_25 = {{3{vector[21]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_22_26 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_26 = {{4{vector[21]}}, vector};
  end
  endfunction


  function automatic [26:0] conv_s2s_22_27 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_27 = {{5{vector[21]}}, vector};
  end
  endfunction


  function automatic [27:0] conv_s2s_22_28 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_28 = {{6{vector[21]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_23_24 ;
    input [22:0]  vector ;
  begin
    conv_s2s_23_24 = {vector[22], vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_23_25 ;
    input [22:0]  vector ;
  begin
    conv_s2s_23_25 = {{2{vector[22]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_23_26 ;
    input [22:0]  vector ;
  begin
    conv_s2s_23_26 = {{3{vector[22]}}, vector};
  end
  endfunction


  function automatic [26:0] conv_s2s_23_27 ;
    input [22:0]  vector ;
  begin
    conv_s2s_23_27 = {{4{vector[22]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_24_25 ;
    input [23:0]  vector ;
  begin
    conv_s2s_24_25 = {vector[23], vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_24_26 ;
    input [23:0]  vector ;
  begin
    conv_s2s_24_26 = {{2{vector[23]}}, vector};
  end
  endfunction


  function automatic [26:0] conv_s2s_24_27 ;
    input [23:0]  vector ;
  begin
    conv_s2s_24_27 = {{3{vector[23]}}, vector};
  end
  endfunction


  function automatic [27:0] conv_s2s_24_28 ;
    input [23:0]  vector ;
  begin
    conv_s2s_24_28 = {{4{vector[23]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_25_26 ;
    input [24:0]  vector ;
  begin
    conv_s2s_25_26 = {vector[24], vector};
  end
  endfunction


  function automatic [27:0] conv_s2s_25_28 ;
    input [24:0]  vector ;
  begin
    conv_s2s_25_28 = {{3{vector[24]}}, vector};
  end
  endfunction


  function automatic [26:0] conv_s2s_26_27 ;
    input [25:0]  vector ;
  begin
    conv_s2s_26_27 = {vector[25], vector};
  end
  endfunction


  function automatic [27:0] conv_s2s_27_28 ;
    input [26:0]  vector ;
  begin
    conv_s2s_27_28 = {vector[26], vector};
  end
  endfunction


  function automatic [8:0] conv_s2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_s2u_8_9 = {vector[7], vector};
  end
  endfunction


  function automatic [9:0] conv_s2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_s2u_9_10 = {vector[8], vector};
  end
  endfunction


  function automatic [10:0] conv_s2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_s2u_10_11 = {vector[9], vector};
  end
  endfunction


  function automatic [11:0] conv_s2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_s2u_11_12 = {vector[10], vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_11_18 ;
    input [10:0]  vector ;
  begin
    conv_s2u_11_18 = {{7{vector[10]}}, vector};
  end
  endfunction


  function automatic [12:0] conv_s2u_12_13 ;
    input [11:0]  vector ;
  begin
    conv_s2u_12_13 = {vector[11], vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_12_18 ;
    input [11:0]  vector ;
  begin
    conv_s2u_12_18 = {{6{vector[11]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_12_19 ;
    input [11:0]  vector ;
  begin
    conv_s2u_12_19 = {{7{vector[11]}}, vector};
  end
  endfunction


  function automatic [13:0] conv_s2u_13_14 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_14 = {vector[12], vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_13_18 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_18 = {{5{vector[12]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_13_19 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_19 = {{6{vector[12]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_14_18 ;
    input [13:0]  vector ;
  begin
    conv_s2u_14_18 = {{4{vector[13]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_14_19 ;
    input [13:0]  vector ;
  begin
    conv_s2u_14_19 = {{5{vector[13]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_15_18 ;
    input [14:0]  vector ;
  begin
    conv_s2u_15_18 = {{3{vector[14]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_15_19 ;
    input [14:0]  vector ;
  begin
    conv_s2u_15_19 = {{4{vector[14]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2u_16_17 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_17 = {vector[15], vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_16_18 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_18 = {{2{vector[15]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_16_19 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_19 = {{3{vector[15]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_17_18 ;
    input [16:0]  vector ;
  begin
    conv_s2u_17_18 = {vector[16], vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_17_19 ;
    input [16:0]  vector ;
  begin
    conv_s2u_17_19 = {{2{vector[16]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_19 = {vector[17], vector};
  end
  endfunction


  function automatic [19:0] conv_s2u_18_20 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_20 = {{2{vector[17]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2u_18_21 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_21 = {{3{vector[17]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_18_22 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_22 = {{4{vector[17]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_18_23 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_23 = {{5{vector[17]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2u_18_24 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_24 = {{6{vector[17]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_18_25 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_25 = {{7{vector[17]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2u_19_20 ;
    input [18:0]  vector ;
  begin
    conv_s2u_19_20 = {vector[18], vector};
  end
  endfunction


  function automatic [20:0] conv_s2u_19_21 ;
    input [18:0]  vector ;
  begin
    conv_s2u_19_21 = {{2{vector[18]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_19_22 ;
    input [18:0]  vector ;
  begin
    conv_s2u_19_22 = {{3{vector[18]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_19_23 ;
    input [18:0]  vector ;
  begin
    conv_s2u_19_23 = {{4{vector[18]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2u_19_24 ;
    input [18:0]  vector ;
  begin
    conv_s2u_19_24 = {{5{vector[18]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2u_20_21 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_21 = {vector[19], vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_20_22 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_22 = {{2{vector[19]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_20_23 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_23 = {{3{vector[19]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2u_20_24 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_24 = {{4{vector[19]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_20_25 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_25 = {{5{vector[19]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_21_22 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_22 = {vector[20], vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_21_23 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_23 = {{2{vector[20]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2u_21_24 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_24 = {{3{vector[20]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2u_21_26 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_26 = {{5{vector[20]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_22_23 ;
    input [21:0]  vector ;
  begin
    conv_s2u_22_23 = {vector[21], vector};
  end
  endfunction


  function automatic [23:0] conv_s2u_22_24 ;
    input [21:0]  vector ;
  begin
    conv_s2u_22_24 = {{2{vector[21]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_22_25 ;
    input [21:0]  vector ;
  begin
    conv_s2u_22_25 = {{3{vector[21]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2u_23_24 ;
    input [22:0]  vector ;
  begin
    conv_s2u_23_24 = {vector[22], vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_23_25 ;
    input [22:0]  vector ;
  begin
    conv_s2u_23_25 = {{2{vector[22]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_24_25 ;
    input [23:0]  vector ;
  begin
    conv_s2u_24_25 = {vector[23], vector};
  end
  endfunction


  function automatic [25:0] conv_s2u_24_26 ;
    input [23:0]  vector ;
  begin
    conv_s2u_24_26 = {{2{vector[23]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2u_25_26 ;
    input [24:0]  vector ;
  begin
    conv_s2u_25_26 = {vector[24], vector};
  end
  endfunction


  function automatic [15:0] conv_u2s_1_16 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_16 = {{15{1'b0}}, vector};
  end
  endfunction


  function automatic [13:0] conv_u2s_11_14 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_14 = {{3{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    nnet_dense_large_input_t_layer2_t_config2
// ------------------------------------------------------------------


module nnet_dense_large_input_t_layer2_t_config2 (
  data_rsc_dat, res_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_srst,
      ccs_ccore_en
);
  input [179:0] data_rsc_dat;
  output [575:0] res_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  nnet_dense_large_input_t_layer2_t_config2_core nnet_dense_large_input_t_layer2_t_config2_core_inst
      (
      .data_rsc_dat(data_rsc_dat),
      .res_rsc_z(res_rsc_z),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4a/835166 Production Release
//  HLS Date:       Thu Sep  5 21:35:46 PDT 2019
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Mon Oct 21 14:04:18 2019
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    keras1layer_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module keras1layer_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [6:0] fsm_output;
  reg [6:0] fsm_output;


  // FSM State Type Declaration for keras1layer_core_core_fsm_1
  parameter
    core_rlp_C_0 = 3'd0,
    main_C_0 = 3'd1,
    main_C_1 = 3'd2,
    main_C_2 = 3'd3,
    main_C_3 = 3'd4,
    main_C_4 = 3'd5,
    main_C_5 = 3'd6;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : keras1layer_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 7'b0000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 7'b0000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 7'b0001000;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 7'b0010000;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 7'b0100000;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 7'b1000000;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 7'b0000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    keras1layer_core_staller
// ------------------------------------------------------------------


module keras1layer_core_staller (
  clk, rst, core_wen, core_wten, input_1_rsci_wen_comp, layer5_out_rsci_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  reg core_wten;
  input input_1_rsci_wen_comp;
  input layer5_out_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = input_1_rsci_wen_comp & layer5_out_rsci_wen_comp;
  always @(posedge clk) begin
    if ( rst ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    keras1layer_core_wait_dp
// ------------------------------------------------------------------


module keras1layer_core_wait_dp (
  ensig_cgo_iro, ensig_cgo_iro_1, ensig_cgo_iro_2, ensig_cgo_iro_3, core_wen, ensig_cgo,
      nnet_sigmoid_layer4_t_result_t_sigmoid_config5_inst_rsci_ccs_ccore_en, ensig_cgo_1,
      nnet_dense_large_layer3_t_layer4_t_config4_cmp_ccs_ccore_en, ensig_cgo_2, nnet_relu_layer2_t_layer3_t_relu_config3_cmp_ccs_ccore_en,
      ensig_cgo_3, nnet_dense_large_input_t_layer2_t_config2_cmp_ccs_ccore_en
);
  input ensig_cgo_iro;
  input ensig_cgo_iro_1;
  input ensig_cgo_iro_2;
  input ensig_cgo_iro_3;
  input core_wen;
  input ensig_cgo;
  output nnet_sigmoid_layer4_t_result_t_sigmoid_config5_inst_rsci_ccs_ccore_en;
  input ensig_cgo_1;
  output nnet_dense_large_layer3_t_layer4_t_config4_cmp_ccs_ccore_en;
  input ensig_cgo_2;
  output nnet_relu_layer2_t_layer3_t_relu_config3_cmp_ccs_ccore_en;
  input ensig_cgo_3;
  output nnet_dense_large_input_t_layer2_t_config2_cmp_ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  assign nnet_sigmoid_layer4_t_result_t_sigmoid_config5_inst_rsci_ccs_ccore_en =
      core_wen & (ensig_cgo | ensig_cgo_iro);
  assign nnet_dense_large_layer3_t_layer4_t_config4_cmp_ccs_ccore_en = core_wen &
      (ensig_cgo_1 | ensig_cgo_iro_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_cmp_ccs_ccore_en = core_wen & (ensig_cgo_2
      | ensig_cgo_iro_2);
  assign nnet_dense_large_input_t_layer2_t_config2_cmp_ccs_ccore_en = core_wen &
      (ensig_cgo_3 | ensig_cgo_iro_3);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    CGHpart
// ------------------------------------------------------------------


module CGHpart (
  CGHpart_isig
);
  input CGHpart_isig;



  // Interconnect Declarations for Component Instantiations 
endmodule

// ------------------------------------------------------------------
//  Design Unit:    keras1layer_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module keras1layer_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl (
  core_wten, const_size_out_1_rsci_iswt0, const_size_out_1_rsci_ivld_core_sct
);
  input core_wten;
  input const_size_out_1_rsci_iswt0;
  output const_size_out_1_rsci_ivld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_out_1_rsci_ivld_core_sct = const_size_out_1_rsci_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    keras1layer_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module keras1layer_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl (
  core_wten, const_size_in_1_rsci_iswt0, const_size_in_1_rsci_ivld_core_sct
);
  input core_wten;
  input const_size_in_1_rsci_iswt0;
  output const_size_in_1_rsci_ivld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_in_1_rsci_ivld_core_sct = const_size_in_1_rsci_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    keras1layer_core_layer5_out_rsci_layer5_out_rsc_wait_dp
// ------------------------------------------------------------------


module keras1layer_core_layer5_out_rsci_layer5_out_rsc_wait_dp (
  clk, rst, layer5_out_rsci_oswt, layer5_out_rsci_wen_comp, layer5_out_rsci_biwt,
      layer5_out_rsci_bdwt, layer5_out_rsci_bcwt
);
  input clk;
  input rst;
  input layer5_out_rsci_oswt;
  output layer5_out_rsci_wen_comp;
  input layer5_out_rsci_biwt;
  input layer5_out_rsci_bdwt;
  output layer5_out_rsci_bcwt;
  reg layer5_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign layer5_out_rsci_wen_comp = (~ layer5_out_rsci_oswt) | layer5_out_rsci_biwt
      | layer5_out_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      layer5_out_rsci_bcwt <= 1'b0;
    end
    else begin
      layer5_out_rsci_bcwt <= ~((~(layer5_out_rsci_bcwt | layer5_out_rsci_biwt))
          | layer5_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    keras1layer_core_layer5_out_rsci_layer5_out_rsc_wait_ctrl
// ------------------------------------------------------------------


module keras1layer_core_layer5_out_rsci_layer5_out_rsc_wait_ctrl (
  core_wen, layer5_out_rsci_oswt, layer5_out_rsci_irdy, layer5_out_rsci_biwt, layer5_out_rsci_bdwt,
      layer5_out_rsci_bcwt, layer5_out_rsci_ivld_core_sct
);
  input core_wen;
  input layer5_out_rsci_oswt;
  input layer5_out_rsci_irdy;
  output layer5_out_rsci_biwt;
  output layer5_out_rsci_bdwt;
  input layer5_out_rsci_bcwt;
  output layer5_out_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire layer5_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign layer5_out_rsci_bdwt = layer5_out_rsci_oswt & core_wen;
  assign layer5_out_rsci_biwt = layer5_out_rsci_ogwt & layer5_out_rsci_irdy;
  assign layer5_out_rsci_ogwt = layer5_out_rsci_oswt & (~ layer5_out_rsci_bcwt);
  assign layer5_out_rsci_ivld_core_sct = layer5_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    keras1layer_core_input_1_rsci_input_1_rsc_wait_dp
// ------------------------------------------------------------------


module keras1layer_core_input_1_rsci_input_1_rsc_wait_dp (
  clk, rst, input_1_rsci_oswt, input_1_rsci_wen_comp, input_1_rsci_idat_mxwt, input_1_rsci_biwt,
      input_1_rsci_bdwt, input_1_rsci_bcwt, input_1_rsci_idat
);
  input clk;
  input rst;
  input input_1_rsci_oswt;
  output input_1_rsci_wen_comp;
  output [179:0] input_1_rsci_idat_mxwt;
  input input_1_rsci_biwt;
  input input_1_rsci_bdwt;
  output input_1_rsci_bcwt;
  reg input_1_rsci_bcwt;
  input [179:0] input_1_rsci_idat;


  // Interconnect Declarations
  reg [179:0] input_1_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_1_rsci_wen_comp = (~ input_1_rsci_oswt) | input_1_rsci_biwt | input_1_rsci_bcwt;
  assign input_1_rsci_idat_mxwt = MUX_v_180_2_2(input_1_rsci_idat, input_1_rsci_idat_bfwt,
      input_1_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      input_1_rsci_bcwt <= 1'b0;
      input_1_rsci_idat_bfwt <= 180'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else begin
      input_1_rsci_bcwt <= ~((~(input_1_rsci_bcwt | input_1_rsci_biwt)) | input_1_rsci_bdwt);
      input_1_rsci_idat_bfwt <= input_1_rsci_idat_mxwt;
    end
  end

  function automatic [179:0] MUX_v_180_2_2;
    input [179:0] input_0;
    input [179:0] input_1;
    input [0:0] sel;
    reg [179:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_180_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    keras1layer_core_input_1_rsci_input_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module keras1layer_core_input_1_rsci_input_1_rsc_wait_ctrl (
  core_wen, input_1_rsci_oswt, input_1_rsci_biwt, input_1_rsci_bdwt, input_1_rsci_bcwt,
      input_1_rsci_irdy_core_sct, input_1_rsci_ivld
);
  input core_wen;
  input input_1_rsci_oswt;
  output input_1_rsci_biwt;
  output input_1_rsci_bdwt;
  input input_1_rsci_bcwt;
  output input_1_rsci_irdy_core_sct;
  input input_1_rsci_ivld;


  // Interconnect Declarations
  wire input_1_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_1_rsci_bdwt = input_1_rsci_oswt & core_wen;
  assign input_1_rsci_biwt = input_1_rsci_ogwt & input_1_rsci_ivld;
  assign input_1_rsci_ogwt = input_1_rsci_oswt & (~ input_1_rsci_bcwt);
  assign input_1_rsci_irdy_core_sct = input_1_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    keras1layer_core_const_size_out_1_rsci
// ------------------------------------------------------------------


module keras1layer_core_const_size_out_1_rsci (
  const_size_out_1_rsc_dat, const_size_out_1_rsc_vld, core_wten, const_size_out_1_rsci_iswt0
);
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  input core_wten;
  input const_size_out_1_rsci_iswt0;


  // Interconnect Declarations
  wire const_size_out_1_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_vld_v1 #(.rscid(32'sd21),
  .width(32'sd16)) const_size_out_1_rsci (
      .ivld(const_size_out_1_rsci_ivld_core_sct),
      .idat(16'b0000000000000001),
      .vld(const_size_out_1_rsc_vld),
      .dat(const_size_out_1_rsc_dat)
    );
  keras1layer_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl keras1layer_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_out_1_rsci_iswt0(const_size_out_1_rsci_iswt0),
      .const_size_out_1_rsci_ivld_core_sct(const_size_out_1_rsci_ivld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    keras1layer_core_const_size_in_1_rsci
// ------------------------------------------------------------------


module keras1layer_core_const_size_in_1_rsci (
  const_size_in_1_rsc_dat, const_size_in_1_rsc_vld, core_wten, const_size_in_1_rsci_iswt0
);
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  input core_wten;
  input const_size_in_1_rsci_iswt0;


  // Interconnect Declarations
  wire const_size_in_1_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_vld_v1 #(.rscid(32'sd20),
  .width(32'sd16)) const_size_in_1_rsci (
      .ivld(const_size_in_1_rsci_ivld_core_sct),
      .idat(16'b0000000000001010),
      .vld(const_size_in_1_rsc_vld),
      .dat(const_size_in_1_rsc_dat)
    );
  keras1layer_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl keras1layer_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_in_1_rsci_iswt0(const_size_in_1_rsci_iswt0),
      .const_size_in_1_rsci_ivld_core_sct(const_size_in_1_rsci_ivld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    keras1layer_core_layer5_out_rsci
// ------------------------------------------------------------------


module keras1layer_core_layer5_out_rsci (
  clk, rst, layer5_out_rsc_dat, layer5_out_rsc_vld, layer5_out_rsc_rdy, core_wen,
      layer5_out_rsci_oswt, layer5_out_rsci_wen_comp, layer5_out_rsci_idat
);
  input clk;
  input rst;
  output [17:0] layer5_out_rsc_dat;
  output layer5_out_rsc_vld;
  input layer5_out_rsc_rdy;
  input core_wen;
  input layer5_out_rsci_oswt;
  output layer5_out_rsci_wen_comp;
  input [17:0] layer5_out_rsci_idat;


  // Interconnect Declarations
  wire layer5_out_rsci_irdy;
  wire layer5_out_rsci_biwt;
  wire layer5_out_rsci_bdwt;
  wire layer5_out_rsci_bcwt;
  wire layer5_out_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd19),
  .width(32'sd18)) layer5_out_rsci (
      .irdy(layer5_out_rsci_irdy),
      .ivld(layer5_out_rsci_ivld_core_sct),
      .idat(layer5_out_rsci_idat),
      .rdy(layer5_out_rsc_rdy),
      .vld(layer5_out_rsc_vld),
      .dat(layer5_out_rsc_dat)
    );
  keras1layer_core_layer5_out_rsci_layer5_out_rsc_wait_ctrl keras1layer_core_layer5_out_rsci_layer5_out_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .layer5_out_rsci_oswt(layer5_out_rsci_oswt),
      .layer5_out_rsci_irdy(layer5_out_rsci_irdy),
      .layer5_out_rsci_biwt(layer5_out_rsci_biwt),
      .layer5_out_rsci_bdwt(layer5_out_rsci_bdwt),
      .layer5_out_rsci_bcwt(layer5_out_rsci_bcwt),
      .layer5_out_rsci_ivld_core_sct(layer5_out_rsci_ivld_core_sct)
    );
  keras1layer_core_layer5_out_rsci_layer5_out_rsc_wait_dp keras1layer_core_layer5_out_rsci_layer5_out_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .layer5_out_rsci_oswt(layer5_out_rsci_oswt),
      .layer5_out_rsci_wen_comp(layer5_out_rsci_wen_comp),
      .layer5_out_rsci_biwt(layer5_out_rsci_biwt),
      .layer5_out_rsci_bdwt(layer5_out_rsci_bdwt),
      .layer5_out_rsci_bcwt(layer5_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    keras1layer_core_input_1_rsci
// ------------------------------------------------------------------


module keras1layer_core_input_1_rsci (
  clk, rst, input_1_rsc_dat, input_1_rsc_vld, input_1_rsc_rdy, core_wen, input_1_rsci_oswt,
      input_1_rsci_wen_comp, input_1_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [179:0] input_1_rsc_dat;
  input input_1_rsc_vld;
  output input_1_rsc_rdy;
  input core_wen;
  input input_1_rsci_oswt;
  output input_1_rsci_wen_comp;
  output [179:0] input_1_rsci_idat_mxwt;


  // Interconnect Declarations
  wire input_1_rsci_biwt;
  wire input_1_rsci_bdwt;
  wire input_1_rsci_bcwt;
  wire input_1_rsci_irdy_core_sct;
  wire input_1_rsci_ivld;
  wire [179:0] input_1_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd18),
  .width(32'sd180)) input_1_rsci (
      .rdy(input_1_rsc_rdy),
      .vld(input_1_rsc_vld),
      .dat(input_1_rsc_dat),
      .irdy(input_1_rsci_irdy_core_sct),
      .ivld(input_1_rsci_ivld),
      .idat(input_1_rsci_idat)
    );
  keras1layer_core_input_1_rsci_input_1_rsc_wait_ctrl keras1layer_core_input_1_rsci_input_1_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .input_1_rsci_oswt(input_1_rsci_oswt),
      .input_1_rsci_biwt(input_1_rsci_biwt),
      .input_1_rsci_bdwt(input_1_rsci_bdwt),
      .input_1_rsci_bcwt(input_1_rsci_bcwt),
      .input_1_rsci_irdy_core_sct(input_1_rsci_irdy_core_sct),
      .input_1_rsci_ivld(input_1_rsci_ivld)
    );
  keras1layer_core_input_1_rsci_input_1_rsc_wait_dp keras1layer_core_input_1_rsci_input_1_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input_1_rsci_oswt(input_1_rsci_oswt),
      .input_1_rsci_wen_comp(input_1_rsci_wen_comp),
      .input_1_rsci_idat_mxwt(input_1_rsci_idat_mxwt),
      .input_1_rsci_biwt(input_1_rsci_biwt),
      .input_1_rsci_bdwt(input_1_rsci_bdwt),
      .input_1_rsci_bcwt(input_1_rsci_bcwt),
      .input_1_rsci_idat(input_1_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    keras1layer_core
// ------------------------------------------------------------------


module keras1layer_core (
  clk, rst, input_1_rsc_dat, input_1_rsc_vld, input_1_rsc_rdy, layer5_out_rsc_dat,
      layer5_out_rsc_vld, layer5_out_rsc_rdy, const_size_in_1_rsc_dat, const_size_in_1_rsc_vld,
      const_size_out_1_rsc_dat, const_size_out_1_rsc_vld
);
  input clk;
  input rst;
  input [179:0] input_1_rsc_dat;
  input input_1_rsc_vld;
  output input_1_rsc_rdy;
  output [17:0] layer5_out_rsc_dat;
  output layer5_out_rsc_vld;
  input layer5_out_rsc_rdy;
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;


  // Interconnect Declarations
  wire core_wen;
  wire core_wten;
  wire input_1_rsci_wen_comp;
  wire [179:0] input_1_rsci_idat_mxwt;
  wire layer5_out_rsci_wen_comp;
  reg [17:0] layer5_out_rsci_idat;
  wire [17:0] nnet_sigmoid_layer4_t_result_t_sigmoid_config5_inst_rsci_res_rsc_z;
  wire nnet_sigmoid_layer4_t_result_t_sigmoid_config5_inst_rsci_ccs_ccore_en;
  wire [17:0] nnet_dense_large_layer3_t_layer4_t_config4_cmp_res_rsc_z;
  wire nnet_dense_large_layer3_t_layer4_t_config4_cmp_ccs_ccore_en;
  wire [575:0] nnet_relu_layer2_t_layer3_t_relu_config3_cmp_res_rsc_z;
  wire nnet_relu_layer2_t_layer3_t_relu_config3_cmp_ccs_ccore_en;
  wire [575:0] nnet_dense_large_input_t_layer2_t_config2_cmp_res_rsc_z;
  wire nnet_dense_large_input_t_layer2_t_config2_cmp_ccs_ccore_en;
  wire [6:0] fsm_output;
  reg reg_const_size_out_1_rsci_ivld_core_psct_cse;
  reg reg_layer5_out_rsci_ivld_core_psct_cse;
  reg reg_ensig_cgo_3_cse;
  reg reg_ensig_cgo_2_cse;
  reg reg_ensig_cgo_1_cse;
  reg reg_ensig_cgo_cse;
  wire or_11_rmff;
  wire or_9_rmff;
  wire or_7_rmff;
  wire or_5_rmff;


  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_nnet_sigmoid_layer4_t_result_t_sigmoid_config5_inst_rsci_ccs_ccore_start_rsc_dat;
  assign nl_nnet_sigmoid_layer4_t_result_t_sigmoid_config5_inst_rsci_ccs_ccore_start_rsc_dat
      = fsm_output[4];
  wire [0:0] nl_nnet_dense_large_layer3_t_layer4_t_config4_cmp_ccs_ccore_start_rsc_dat;
  assign nl_nnet_dense_large_layer3_t_layer4_t_config4_cmp_ccs_ccore_start_rsc_dat
      = fsm_output[3];
  wire [0:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_cmp_ccs_ccore_start_rsc_dat;
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_cmp_ccs_ccore_start_rsc_dat
      = fsm_output[2];
  wire [0:0] nl_nnet_dense_large_input_t_layer2_t_config2_cmp_ccs_ccore_start_rsc_dat;
  assign nl_nnet_dense_large_input_t_layer2_t_config2_cmp_ccs_ccore_start_rsc_dat
      = fsm_output[1];
  nnet_sigmoid_layer4_t_result_t_sigmoid_config5  nnet_sigmoid_layer4_t_result_t_sigmoid_config5_inst_rsci
      (
      .data_rsc_dat(nnet_dense_large_layer3_t_layer4_t_config4_cmp_res_rsc_z),
      .res_rsc_z(nnet_sigmoid_layer4_t_result_t_sigmoid_config5_inst_rsci_res_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(nnet_sigmoid_layer4_t_result_t_sigmoid_config5_inst_rsci_ccs_ccore_en),
      .ccs_ccore_srst(rst),
      .ccs_ccore_start_rsc_dat(nl_nnet_sigmoid_layer4_t_result_t_sigmoid_config5_inst_rsci_ccs_ccore_start_rsc_dat[0:0])
    );
  nnet_dense_large_layer3_t_layer4_t_config4  nnet_dense_large_layer3_t_layer4_t_config4_cmp
      (
      .data_rsc_dat(nnet_relu_layer2_t_layer3_t_relu_config3_cmp_res_rsc_z),
      .res_rsc_z(nnet_dense_large_layer3_t_layer4_t_config4_cmp_res_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(nnet_dense_large_layer3_t_layer4_t_config4_cmp_ccs_ccore_en),
      .ccs_ccore_srst(rst),
      .ccs_ccore_start_rsc_dat(nl_nnet_dense_large_layer3_t_layer4_t_config4_cmp_ccs_ccore_start_rsc_dat[0:0])
    );
  nnet_relu_layer2_t_layer3_t_relu_config3  nnet_relu_layer2_t_layer3_t_relu_config3_cmp
      (
      .data_rsc_dat(nnet_dense_large_input_t_layer2_t_config2_cmp_res_rsc_z),
      .res_rsc_z(nnet_relu_layer2_t_layer3_t_relu_config3_cmp_res_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(nnet_relu_layer2_t_layer3_t_relu_config3_cmp_ccs_ccore_en),
      .ccs_ccore_srst(rst),
      .ccs_ccore_start_rsc_dat(nl_nnet_relu_layer2_t_layer3_t_relu_config3_cmp_ccs_ccore_start_rsc_dat[0:0])
    );
  nnet_dense_large_input_t_layer2_t_config2  nnet_dense_large_input_t_layer2_t_config2_cmp
      (
      .data_rsc_dat(input_1_rsci_idat_mxwt),
      .res_rsc_z(nnet_dense_large_input_t_layer2_t_config2_cmp_res_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(nnet_dense_large_input_t_layer2_t_config2_cmp_ccs_ccore_en),
      .ccs_ccore_srst(rst),
      .ccs_ccore_start_rsc_dat(nl_nnet_dense_large_input_t_layer2_t_config2_cmp_ccs_ccore_start_rsc_dat[0:0])
    );
  keras1layer_core_input_1_rsci keras1layer_core_input_1_rsci_inst (
      .clk(clk),
      .rst(rst),
      .input_1_rsc_dat(input_1_rsc_dat),
      .input_1_rsc_vld(input_1_rsc_vld),
      .input_1_rsc_rdy(input_1_rsc_rdy),
      .core_wen(core_wen),
      .input_1_rsci_oswt(reg_const_size_out_1_rsci_ivld_core_psct_cse),
      .input_1_rsci_wen_comp(input_1_rsci_wen_comp),
      .input_1_rsci_idat_mxwt(input_1_rsci_idat_mxwt)
    );
  keras1layer_core_layer5_out_rsci keras1layer_core_layer5_out_rsci_inst (
      .clk(clk),
      .rst(rst),
      .layer5_out_rsc_dat(layer5_out_rsc_dat),
      .layer5_out_rsc_vld(layer5_out_rsc_vld),
      .layer5_out_rsc_rdy(layer5_out_rsc_rdy),
      .core_wen(core_wen),
      .layer5_out_rsci_oswt(reg_layer5_out_rsci_ivld_core_psct_cse),
      .layer5_out_rsci_wen_comp(layer5_out_rsci_wen_comp),
      .layer5_out_rsci_idat(layer5_out_rsci_idat)
    );
  keras1layer_core_const_size_in_1_rsci keras1layer_core_const_size_in_1_rsci_inst
      (
      .const_size_in_1_rsc_dat(const_size_in_1_rsc_dat),
      .const_size_in_1_rsc_vld(const_size_in_1_rsc_vld),
      .core_wten(core_wten),
      .const_size_in_1_rsci_iswt0(reg_const_size_out_1_rsci_ivld_core_psct_cse)
    );
  keras1layer_core_const_size_out_1_rsci keras1layer_core_const_size_out_1_rsci_inst
      (
      .const_size_out_1_rsc_dat(const_size_out_1_rsc_dat),
      .const_size_out_1_rsc_vld(const_size_out_1_rsc_vld),
      .core_wten(core_wten),
      .const_size_out_1_rsci_iswt0(reg_const_size_out_1_rsci_ivld_core_psct_cse)
    );
  keras1layer_core_wait_dp keras1layer_core_wait_dp_inst (
      .ensig_cgo_iro(or_11_rmff),
      .ensig_cgo_iro_1(or_9_rmff),
      .ensig_cgo_iro_2(or_7_rmff),
      .ensig_cgo_iro_3(or_5_rmff),
      .core_wen(core_wen),
      .ensig_cgo(reg_ensig_cgo_cse),
      .nnet_sigmoid_layer4_t_result_t_sigmoid_config5_inst_rsci_ccs_ccore_en(nnet_sigmoid_layer4_t_result_t_sigmoid_config5_inst_rsci_ccs_ccore_en),
      .ensig_cgo_1(reg_ensig_cgo_1_cse),
      .nnet_dense_large_layer3_t_layer4_t_config4_cmp_ccs_ccore_en(nnet_dense_large_layer3_t_layer4_t_config4_cmp_ccs_ccore_en),
      .ensig_cgo_2(reg_ensig_cgo_2_cse),
      .nnet_relu_layer2_t_layer3_t_relu_config3_cmp_ccs_ccore_en(nnet_relu_layer2_t_layer3_t_relu_config3_cmp_ccs_ccore_en),
      .ensig_cgo_3(reg_ensig_cgo_3_cse),
      .nnet_dense_large_input_t_layer2_t_config2_cmp_ccs_ccore_en(nnet_dense_large_input_t_layer2_t_config2_cmp_ccs_ccore_en)
    );
  keras1layer_core_staller keras1layer_core_staller_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .input_1_rsci_wen_comp(input_1_rsci_wen_comp),
      .layer5_out_rsci_wen_comp(layer5_out_rsci_wen_comp)
    );
  keras1layer_core_core_fsm keras1layer_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign or_5_rmff = (fsm_output[2:1]!=2'b00);
  assign or_7_rmff = (fsm_output[3:2]!=2'b00);
  assign or_9_rmff = (fsm_output[4:3]!=2'b00);
  assign or_11_rmff = (fsm_output[5:4]!=2'b00);
  always @(posedge clk) begin
    if ( rst ) begin
      reg_ensig_cgo_3_cse <= 1'b0;
      reg_ensig_cgo_2_cse <= 1'b0;
      reg_ensig_cgo_1_cse <= 1'b0;
      reg_ensig_cgo_cse <= 1'b0;
      reg_const_size_out_1_rsci_ivld_core_psct_cse <= 1'b0;
      reg_layer5_out_rsci_ivld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_ensig_cgo_3_cse <= or_5_rmff;
      reg_ensig_cgo_2_cse <= or_7_rmff;
      reg_ensig_cgo_1_cse <= or_9_rmff;
      reg_ensig_cgo_cse <= or_11_rmff;
      reg_const_size_out_1_rsci_ivld_core_psct_cse <= (fsm_output[6]) | (fsm_output[0]);
      reg_layer5_out_rsci_ivld_core_psct_cse <= fsm_output[5];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer5_out_rsci_idat <= 18'b000000000000000000;
    end
    else if ( core_wen & (fsm_output[5]) ) begin
      layer5_out_rsci_idat <= nnet_sigmoid_layer4_t_result_t_sigmoid_config5_inst_rsci_res_rsc_z;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    keras1layer
// ------------------------------------------------------------------


module keras1layer (
  clk, rst, input_1_rsc_dat, input_1_rsc_vld, input_1_rsc_rdy, layer5_out_rsc_dat,
      layer5_out_rsc_vld, layer5_out_rsc_rdy, const_size_in_1_rsc_dat, const_size_in_1_rsc_vld,
      const_size_out_1_rsc_dat, const_size_out_1_rsc_vld
);
  input clk;
  input rst;
  input [179:0] input_1_rsc_dat;
  input input_1_rsc_vld;
  output input_1_rsc_rdy;
  output [17:0] layer5_out_rsc_dat;
  output layer5_out_rsc_vld;
  input layer5_out_rsc_rdy;
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;



  // Interconnect Declarations for Component Instantiations 
  keras1layer_core keras1layer_core_inst (
      .clk(clk),
      .rst(rst),
      .input_1_rsc_dat(input_1_rsc_dat),
      .input_1_rsc_vld(input_1_rsc_vld),
      .input_1_rsc_rdy(input_1_rsc_rdy),
      .layer5_out_rsc_dat(layer5_out_rsc_dat),
      .layer5_out_rsc_vld(layer5_out_rsc_vld),
      .layer5_out_rsc_rdy(layer5_out_rsc_rdy),
      .const_size_in_1_rsc_dat(const_size_in_1_rsc_dat),
      .const_size_in_1_rsc_vld(const_size_in_1_rsc_vld),
      .const_size_out_1_rsc_dat(const_size_out_1_rsc_dat),
      .const_size_out_1_rsc_vld(const_size_out_1_rsc_vld)
    );
endmodule



