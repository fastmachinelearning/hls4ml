
//------> /opt/cad/catapult/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> /opt/cad/catapult/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  assign dat = idat;
  assign irdy = rdy;
  assign vld = ivld;

endmodule



//------> /opt/cad/catapult/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ../td_ccore_solutions/ROM_1i3_1o10_2c1f806487d17904bea969f4e53173bcb1_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Fri Nov  1 23:14:12 2019
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i3_1o10_2c1f806487d17904bea969f4e53173bcb1
// ------------------------------------------------------------------


module ROM_1i3_1o10_2c1f806487d17904bea969f4e53173bcb1 (
  I_1, O_1
);
  input [2:0] I_1;
  output [9:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_10_8_2(10'b1111111101, 10'b1100011001, 10'b1001100100, 10'b0111010000,
      10'b0101010100, 10'b0011101011, 10'b0010010001, 10'b0001000100, I_1);

  function automatic [9:0] MUX_v_10_8_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [9:0] input_2;
    input [9:0] input_3;
    input [9:0] input_4;
    input [9:0] input_5;
    input [9:0] input_6;
    input [9:0] input_7;
    input [2:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_10_8_2 = result;
  end
  endfunction

endmodule




//------> /opt/cad/catapult/pkgs/siflibs/mgc_shift_br_beh_v5.v 
module mgc_shift_br_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_s(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_s(a,s,1'b0);
     end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshr_u

   //Shift right - signed shift argument
   function [width_z-1:0] fshr_s;
     input [width_a-1:0] arg1;
     input [width_s-1:0] arg2;
     input sbit;
     begin
       if ( arg2[width_s-1] == 1'b0 )
       begin
         fshr_s = fshr_u(arg1, arg2, sbit);
       end
       else
       begin
         fshr_s = fshl_u_1({arg1, 1'b0},~arg2, sbit);
       end
     end
   endfunction 

endmodule

//------> ../td_ccore_solutions/ROM_1i11_1o5_35e12f400da6925eda56234f89e8055db3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Sat Nov  2 10:28:43 2019
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i11_1o5_35e12f400da6925eda56234f89e8055db3
// ------------------------------------------------------------------


module ROM_1i11_1o5_35e12f400da6925eda56234f89e8055db3 (
  I_1, O_1
);
  input [10:0] I_1;
  output [4:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_5_2048_2(5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000,
      5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000,
      5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000,
      5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000,
      5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000,
      5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000,
      5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000,
      5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000,
      5'b00000, 5'b00000, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001,
      5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001,
      5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001,
      5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001,
      5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001,
      5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001,
      5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001,
      5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001,
      5'b00001, 5'b00001, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010,
      5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010,
      5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010,
      5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010,
      5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010,
      5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010,
      5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010,
      5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010,
      5'b00010, 5'b00010, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011,
      5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011,
      5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011,
      5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011,
      5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011,
      5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011,
      5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011,
      5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011,
      5'b00011, 5'b00011, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100,
      5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100,
      5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100,
      5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100,
      5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100,
      5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100,
      5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100,
      5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100,
      5'b00100, 5'b00100, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101,
      5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101,
      5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101,
      5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101,
      5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101,
      5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101,
      5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101,
      5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101,
      5'b00101, 5'b00101, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110,
      5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110,
      5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110,
      5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110,
      5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110,
      5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110,
      5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110,
      5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110,
      5'b00110, 5'b00110, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111,
      5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111,
      5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111,
      5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111,
      5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111,
      5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111,
      5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111,
      5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00111,
      5'b00111, 5'b00111, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000,
      5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000,
      5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000,
      5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000,
      5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000,
      5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000,
      5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000,
      5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b01000,
      5'b01000, 5'b01000, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001,
      5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001,
      5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001,
      5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001,
      5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001,
      5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001,
      5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001,
      5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001,
      5'b01001, 5'b01001, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010,
      5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010,
      5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010,
      5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010,
      5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010,
      5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010,
      5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010,
      5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01010,
      5'b01010, 5'b01010, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011,
      5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011,
      5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011,
      5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011,
      5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011,
      5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011,
      5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011,
      5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011,
      5'b01011, 5'b01011, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100,
      5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100,
      5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100,
      5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100,
      5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100,
      5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100,
      5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100,
      5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01100,
      5'b01100, 5'b01100, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101,
      5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101,
      5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101,
      5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101,
      5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101,
      5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101,
      5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101,
      5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101,
      5'b01101, 5'b01101, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110,
      5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110,
      5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110,
      5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110,
      5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110,
      5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110,
      5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110,
      5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110,
      5'b01110, 5'b01110, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111,
      5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111,
      5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111,
      5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111,
      5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111,
      5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111,
      5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111,
      5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b01111,
      5'b01111, 5'b01111, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000,
      5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000,
      5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000,
      5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000,
      5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000,
      5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000,
      5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000,
      5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000,
      5'b10000, 5'b10000, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001,
      5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001,
      5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001,
      5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001,
      5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001,
      5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001,
      5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001,
      5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001,
      5'b10001, 5'b10001, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010,
      5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010,
      5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010,
      5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010,
      5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010,
      5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010,
      5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010,
      5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b10010,
      5'b10010, 5'b10010, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011,
      5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011,
      5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011,
      5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011,
      5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011,
      5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011,
      5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011,
      5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10011,
      5'b10011, 5'b10011, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100,
      5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100,
      5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100,
      5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100,
      5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100,
      5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100,
      5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100,
      5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100, 5'b10100,
      5'b10100, 5'b10100, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101,
      5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101,
      5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101,
      5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101,
      5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101,
      5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101,
      5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101,
      5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10101,
      5'b10101, 5'b10101, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110,
      5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110,
      5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110,
      5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110,
      5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110,
      5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110,
      5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110,
      5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110,
      5'b10110, 5'b10110, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111,
      5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111,
      5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111,
      5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111,
      5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111,
      5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111,
      5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111,
      5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111, 5'b10111,
      5'b10111, 5'b10111, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000,
      5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000,
      5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000,
      5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000,
      5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000,
      5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000,
      5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000,
      5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000, 5'b11000,
      5'b11000, 5'b11000, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001,
      5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001,
      5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001,
      5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001,
      5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001,
      5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001,
      5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001,
      5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001, 5'b11001,
      5'b11001, 5'b11001, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010,
      5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010,
      5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010,
      5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010,
      5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010,
      5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010,
      5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010,
      5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010, 5'b11010,
      5'b11010, 5'b11010, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011,
      5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011,
      5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011,
      5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011,
      5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011,
      5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011,
      5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011,
      5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011, 5'b11011,
      5'b11011, 5'b11011, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100,
      5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100,
      5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100,
      5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100,
      5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100,
      5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100,
      5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100,
      5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100, 5'b11100,
      5'b11100, 5'b11100, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101,
      5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101,
      5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101,
      5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101,
      5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101,
      5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101,
      5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101,
      5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101, 5'b11101,
      5'b11101, 5'b11101, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110,
      5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110,
      5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110,
      5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110,
      5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110,
      5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110,
      5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110,
      5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110, 5'b11110,
      5'b11110, 5'b11110, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111,
      5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111,
      5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111,
      5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111,
      5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111,
      5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111,
      5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111,
      5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111, 5'b11111,
      5'b11111, 5'b11111, I_1);

  function automatic [4:0] MUX_v_5_2048_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [4:0] input_2;
    input [4:0] input_3;
    input [4:0] input_4;
    input [4:0] input_5;
    input [4:0] input_6;
    input [4:0] input_7;
    input [4:0] input_8;
    input [4:0] input_9;
    input [4:0] input_10;
    input [4:0] input_11;
    input [4:0] input_12;
    input [4:0] input_13;
    input [4:0] input_14;
    input [4:0] input_15;
    input [4:0] input_16;
    input [4:0] input_17;
    input [4:0] input_18;
    input [4:0] input_19;
    input [4:0] input_20;
    input [4:0] input_21;
    input [4:0] input_22;
    input [4:0] input_23;
    input [4:0] input_24;
    input [4:0] input_25;
    input [4:0] input_26;
    input [4:0] input_27;
    input [4:0] input_28;
    input [4:0] input_29;
    input [4:0] input_30;
    input [4:0] input_31;
    input [4:0] input_32;
    input [4:0] input_33;
    input [4:0] input_34;
    input [4:0] input_35;
    input [4:0] input_36;
    input [4:0] input_37;
    input [4:0] input_38;
    input [4:0] input_39;
    input [4:0] input_40;
    input [4:0] input_41;
    input [4:0] input_42;
    input [4:0] input_43;
    input [4:0] input_44;
    input [4:0] input_45;
    input [4:0] input_46;
    input [4:0] input_47;
    input [4:0] input_48;
    input [4:0] input_49;
    input [4:0] input_50;
    input [4:0] input_51;
    input [4:0] input_52;
    input [4:0] input_53;
    input [4:0] input_54;
    input [4:0] input_55;
    input [4:0] input_56;
    input [4:0] input_57;
    input [4:0] input_58;
    input [4:0] input_59;
    input [4:0] input_60;
    input [4:0] input_61;
    input [4:0] input_62;
    input [4:0] input_63;
    input [4:0] input_64;
    input [4:0] input_65;
    input [4:0] input_66;
    input [4:0] input_67;
    input [4:0] input_68;
    input [4:0] input_69;
    input [4:0] input_70;
    input [4:0] input_71;
    input [4:0] input_72;
    input [4:0] input_73;
    input [4:0] input_74;
    input [4:0] input_75;
    input [4:0] input_76;
    input [4:0] input_77;
    input [4:0] input_78;
    input [4:0] input_79;
    input [4:0] input_80;
    input [4:0] input_81;
    input [4:0] input_82;
    input [4:0] input_83;
    input [4:0] input_84;
    input [4:0] input_85;
    input [4:0] input_86;
    input [4:0] input_87;
    input [4:0] input_88;
    input [4:0] input_89;
    input [4:0] input_90;
    input [4:0] input_91;
    input [4:0] input_92;
    input [4:0] input_93;
    input [4:0] input_94;
    input [4:0] input_95;
    input [4:0] input_96;
    input [4:0] input_97;
    input [4:0] input_98;
    input [4:0] input_99;
    input [4:0] input_100;
    input [4:0] input_101;
    input [4:0] input_102;
    input [4:0] input_103;
    input [4:0] input_104;
    input [4:0] input_105;
    input [4:0] input_106;
    input [4:0] input_107;
    input [4:0] input_108;
    input [4:0] input_109;
    input [4:0] input_110;
    input [4:0] input_111;
    input [4:0] input_112;
    input [4:0] input_113;
    input [4:0] input_114;
    input [4:0] input_115;
    input [4:0] input_116;
    input [4:0] input_117;
    input [4:0] input_118;
    input [4:0] input_119;
    input [4:0] input_120;
    input [4:0] input_121;
    input [4:0] input_122;
    input [4:0] input_123;
    input [4:0] input_124;
    input [4:0] input_125;
    input [4:0] input_126;
    input [4:0] input_127;
    input [4:0] input_128;
    input [4:0] input_129;
    input [4:0] input_130;
    input [4:0] input_131;
    input [4:0] input_132;
    input [4:0] input_133;
    input [4:0] input_134;
    input [4:0] input_135;
    input [4:0] input_136;
    input [4:0] input_137;
    input [4:0] input_138;
    input [4:0] input_139;
    input [4:0] input_140;
    input [4:0] input_141;
    input [4:0] input_142;
    input [4:0] input_143;
    input [4:0] input_144;
    input [4:0] input_145;
    input [4:0] input_146;
    input [4:0] input_147;
    input [4:0] input_148;
    input [4:0] input_149;
    input [4:0] input_150;
    input [4:0] input_151;
    input [4:0] input_152;
    input [4:0] input_153;
    input [4:0] input_154;
    input [4:0] input_155;
    input [4:0] input_156;
    input [4:0] input_157;
    input [4:0] input_158;
    input [4:0] input_159;
    input [4:0] input_160;
    input [4:0] input_161;
    input [4:0] input_162;
    input [4:0] input_163;
    input [4:0] input_164;
    input [4:0] input_165;
    input [4:0] input_166;
    input [4:0] input_167;
    input [4:0] input_168;
    input [4:0] input_169;
    input [4:0] input_170;
    input [4:0] input_171;
    input [4:0] input_172;
    input [4:0] input_173;
    input [4:0] input_174;
    input [4:0] input_175;
    input [4:0] input_176;
    input [4:0] input_177;
    input [4:0] input_178;
    input [4:0] input_179;
    input [4:0] input_180;
    input [4:0] input_181;
    input [4:0] input_182;
    input [4:0] input_183;
    input [4:0] input_184;
    input [4:0] input_185;
    input [4:0] input_186;
    input [4:0] input_187;
    input [4:0] input_188;
    input [4:0] input_189;
    input [4:0] input_190;
    input [4:0] input_191;
    input [4:0] input_192;
    input [4:0] input_193;
    input [4:0] input_194;
    input [4:0] input_195;
    input [4:0] input_196;
    input [4:0] input_197;
    input [4:0] input_198;
    input [4:0] input_199;
    input [4:0] input_200;
    input [4:0] input_201;
    input [4:0] input_202;
    input [4:0] input_203;
    input [4:0] input_204;
    input [4:0] input_205;
    input [4:0] input_206;
    input [4:0] input_207;
    input [4:0] input_208;
    input [4:0] input_209;
    input [4:0] input_210;
    input [4:0] input_211;
    input [4:0] input_212;
    input [4:0] input_213;
    input [4:0] input_214;
    input [4:0] input_215;
    input [4:0] input_216;
    input [4:0] input_217;
    input [4:0] input_218;
    input [4:0] input_219;
    input [4:0] input_220;
    input [4:0] input_221;
    input [4:0] input_222;
    input [4:0] input_223;
    input [4:0] input_224;
    input [4:0] input_225;
    input [4:0] input_226;
    input [4:0] input_227;
    input [4:0] input_228;
    input [4:0] input_229;
    input [4:0] input_230;
    input [4:0] input_231;
    input [4:0] input_232;
    input [4:0] input_233;
    input [4:0] input_234;
    input [4:0] input_235;
    input [4:0] input_236;
    input [4:0] input_237;
    input [4:0] input_238;
    input [4:0] input_239;
    input [4:0] input_240;
    input [4:0] input_241;
    input [4:0] input_242;
    input [4:0] input_243;
    input [4:0] input_244;
    input [4:0] input_245;
    input [4:0] input_246;
    input [4:0] input_247;
    input [4:0] input_248;
    input [4:0] input_249;
    input [4:0] input_250;
    input [4:0] input_251;
    input [4:0] input_252;
    input [4:0] input_253;
    input [4:0] input_254;
    input [4:0] input_255;
    input [4:0] input_256;
    input [4:0] input_257;
    input [4:0] input_258;
    input [4:0] input_259;
    input [4:0] input_260;
    input [4:0] input_261;
    input [4:0] input_262;
    input [4:0] input_263;
    input [4:0] input_264;
    input [4:0] input_265;
    input [4:0] input_266;
    input [4:0] input_267;
    input [4:0] input_268;
    input [4:0] input_269;
    input [4:0] input_270;
    input [4:0] input_271;
    input [4:0] input_272;
    input [4:0] input_273;
    input [4:0] input_274;
    input [4:0] input_275;
    input [4:0] input_276;
    input [4:0] input_277;
    input [4:0] input_278;
    input [4:0] input_279;
    input [4:0] input_280;
    input [4:0] input_281;
    input [4:0] input_282;
    input [4:0] input_283;
    input [4:0] input_284;
    input [4:0] input_285;
    input [4:0] input_286;
    input [4:0] input_287;
    input [4:0] input_288;
    input [4:0] input_289;
    input [4:0] input_290;
    input [4:0] input_291;
    input [4:0] input_292;
    input [4:0] input_293;
    input [4:0] input_294;
    input [4:0] input_295;
    input [4:0] input_296;
    input [4:0] input_297;
    input [4:0] input_298;
    input [4:0] input_299;
    input [4:0] input_300;
    input [4:0] input_301;
    input [4:0] input_302;
    input [4:0] input_303;
    input [4:0] input_304;
    input [4:0] input_305;
    input [4:0] input_306;
    input [4:0] input_307;
    input [4:0] input_308;
    input [4:0] input_309;
    input [4:0] input_310;
    input [4:0] input_311;
    input [4:0] input_312;
    input [4:0] input_313;
    input [4:0] input_314;
    input [4:0] input_315;
    input [4:0] input_316;
    input [4:0] input_317;
    input [4:0] input_318;
    input [4:0] input_319;
    input [4:0] input_320;
    input [4:0] input_321;
    input [4:0] input_322;
    input [4:0] input_323;
    input [4:0] input_324;
    input [4:0] input_325;
    input [4:0] input_326;
    input [4:0] input_327;
    input [4:0] input_328;
    input [4:0] input_329;
    input [4:0] input_330;
    input [4:0] input_331;
    input [4:0] input_332;
    input [4:0] input_333;
    input [4:0] input_334;
    input [4:0] input_335;
    input [4:0] input_336;
    input [4:0] input_337;
    input [4:0] input_338;
    input [4:0] input_339;
    input [4:0] input_340;
    input [4:0] input_341;
    input [4:0] input_342;
    input [4:0] input_343;
    input [4:0] input_344;
    input [4:0] input_345;
    input [4:0] input_346;
    input [4:0] input_347;
    input [4:0] input_348;
    input [4:0] input_349;
    input [4:0] input_350;
    input [4:0] input_351;
    input [4:0] input_352;
    input [4:0] input_353;
    input [4:0] input_354;
    input [4:0] input_355;
    input [4:0] input_356;
    input [4:0] input_357;
    input [4:0] input_358;
    input [4:0] input_359;
    input [4:0] input_360;
    input [4:0] input_361;
    input [4:0] input_362;
    input [4:0] input_363;
    input [4:0] input_364;
    input [4:0] input_365;
    input [4:0] input_366;
    input [4:0] input_367;
    input [4:0] input_368;
    input [4:0] input_369;
    input [4:0] input_370;
    input [4:0] input_371;
    input [4:0] input_372;
    input [4:0] input_373;
    input [4:0] input_374;
    input [4:0] input_375;
    input [4:0] input_376;
    input [4:0] input_377;
    input [4:0] input_378;
    input [4:0] input_379;
    input [4:0] input_380;
    input [4:0] input_381;
    input [4:0] input_382;
    input [4:0] input_383;
    input [4:0] input_384;
    input [4:0] input_385;
    input [4:0] input_386;
    input [4:0] input_387;
    input [4:0] input_388;
    input [4:0] input_389;
    input [4:0] input_390;
    input [4:0] input_391;
    input [4:0] input_392;
    input [4:0] input_393;
    input [4:0] input_394;
    input [4:0] input_395;
    input [4:0] input_396;
    input [4:0] input_397;
    input [4:0] input_398;
    input [4:0] input_399;
    input [4:0] input_400;
    input [4:0] input_401;
    input [4:0] input_402;
    input [4:0] input_403;
    input [4:0] input_404;
    input [4:0] input_405;
    input [4:0] input_406;
    input [4:0] input_407;
    input [4:0] input_408;
    input [4:0] input_409;
    input [4:0] input_410;
    input [4:0] input_411;
    input [4:0] input_412;
    input [4:0] input_413;
    input [4:0] input_414;
    input [4:0] input_415;
    input [4:0] input_416;
    input [4:0] input_417;
    input [4:0] input_418;
    input [4:0] input_419;
    input [4:0] input_420;
    input [4:0] input_421;
    input [4:0] input_422;
    input [4:0] input_423;
    input [4:0] input_424;
    input [4:0] input_425;
    input [4:0] input_426;
    input [4:0] input_427;
    input [4:0] input_428;
    input [4:0] input_429;
    input [4:0] input_430;
    input [4:0] input_431;
    input [4:0] input_432;
    input [4:0] input_433;
    input [4:0] input_434;
    input [4:0] input_435;
    input [4:0] input_436;
    input [4:0] input_437;
    input [4:0] input_438;
    input [4:0] input_439;
    input [4:0] input_440;
    input [4:0] input_441;
    input [4:0] input_442;
    input [4:0] input_443;
    input [4:0] input_444;
    input [4:0] input_445;
    input [4:0] input_446;
    input [4:0] input_447;
    input [4:0] input_448;
    input [4:0] input_449;
    input [4:0] input_450;
    input [4:0] input_451;
    input [4:0] input_452;
    input [4:0] input_453;
    input [4:0] input_454;
    input [4:0] input_455;
    input [4:0] input_456;
    input [4:0] input_457;
    input [4:0] input_458;
    input [4:0] input_459;
    input [4:0] input_460;
    input [4:0] input_461;
    input [4:0] input_462;
    input [4:0] input_463;
    input [4:0] input_464;
    input [4:0] input_465;
    input [4:0] input_466;
    input [4:0] input_467;
    input [4:0] input_468;
    input [4:0] input_469;
    input [4:0] input_470;
    input [4:0] input_471;
    input [4:0] input_472;
    input [4:0] input_473;
    input [4:0] input_474;
    input [4:0] input_475;
    input [4:0] input_476;
    input [4:0] input_477;
    input [4:0] input_478;
    input [4:0] input_479;
    input [4:0] input_480;
    input [4:0] input_481;
    input [4:0] input_482;
    input [4:0] input_483;
    input [4:0] input_484;
    input [4:0] input_485;
    input [4:0] input_486;
    input [4:0] input_487;
    input [4:0] input_488;
    input [4:0] input_489;
    input [4:0] input_490;
    input [4:0] input_491;
    input [4:0] input_492;
    input [4:0] input_493;
    input [4:0] input_494;
    input [4:0] input_495;
    input [4:0] input_496;
    input [4:0] input_497;
    input [4:0] input_498;
    input [4:0] input_499;
    input [4:0] input_500;
    input [4:0] input_501;
    input [4:0] input_502;
    input [4:0] input_503;
    input [4:0] input_504;
    input [4:0] input_505;
    input [4:0] input_506;
    input [4:0] input_507;
    input [4:0] input_508;
    input [4:0] input_509;
    input [4:0] input_510;
    input [4:0] input_511;
    input [4:0] input_512;
    input [4:0] input_513;
    input [4:0] input_514;
    input [4:0] input_515;
    input [4:0] input_516;
    input [4:0] input_517;
    input [4:0] input_518;
    input [4:0] input_519;
    input [4:0] input_520;
    input [4:0] input_521;
    input [4:0] input_522;
    input [4:0] input_523;
    input [4:0] input_524;
    input [4:0] input_525;
    input [4:0] input_526;
    input [4:0] input_527;
    input [4:0] input_528;
    input [4:0] input_529;
    input [4:0] input_530;
    input [4:0] input_531;
    input [4:0] input_532;
    input [4:0] input_533;
    input [4:0] input_534;
    input [4:0] input_535;
    input [4:0] input_536;
    input [4:0] input_537;
    input [4:0] input_538;
    input [4:0] input_539;
    input [4:0] input_540;
    input [4:0] input_541;
    input [4:0] input_542;
    input [4:0] input_543;
    input [4:0] input_544;
    input [4:0] input_545;
    input [4:0] input_546;
    input [4:0] input_547;
    input [4:0] input_548;
    input [4:0] input_549;
    input [4:0] input_550;
    input [4:0] input_551;
    input [4:0] input_552;
    input [4:0] input_553;
    input [4:0] input_554;
    input [4:0] input_555;
    input [4:0] input_556;
    input [4:0] input_557;
    input [4:0] input_558;
    input [4:0] input_559;
    input [4:0] input_560;
    input [4:0] input_561;
    input [4:0] input_562;
    input [4:0] input_563;
    input [4:0] input_564;
    input [4:0] input_565;
    input [4:0] input_566;
    input [4:0] input_567;
    input [4:0] input_568;
    input [4:0] input_569;
    input [4:0] input_570;
    input [4:0] input_571;
    input [4:0] input_572;
    input [4:0] input_573;
    input [4:0] input_574;
    input [4:0] input_575;
    input [4:0] input_576;
    input [4:0] input_577;
    input [4:0] input_578;
    input [4:0] input_579;
    input [4:0] input_580;
    input [4:0] input_581;
    input [4:0] input_582;
    input [4:0] input_583;
    input [4:0] input_584;
    input [4:0] input_585;
    input [4:0] input_586;
    input [4:0] input_587;
    input [4:0] input_588;
    input [4:0] input_589;
    input [4:0] input_590;
    input [4:0] input_591;
    input [4:0] input_592;
    input [4:0] input_593;
    input [4:0] input_594;
    input [4:0] input_595;
    input [4:0] input_596;
    input [4:0] input_597;
    input [4:0] input_598;
    input [4:0] input_599;
    input [4:0] input_600;
    input [4:0] input_601;
    input [4:0] input_602;
    input [4:0] input_603;
    input [4:0] input_604;
    input [4:0] input_605;
    input [4:0] input_606;
    input [4:0] input_607;
    input [4:0] input_608;
    input [4:0] input_609;
    input [4:0] input_610;
    input [4:0] input_611;
    input [4:0] input_612;
    input [4:0] input_613;
    input [4:0] input_614;
    input [4:0] input_615;
    input [4:0] input_616;
    input [4:0] input_617;
    input [4:0] input_618;
    input [4:0] input_619;
    input [4:0] input_620;
    input [4:0] input_621;
    input [4:0] input_622;
    input [4:0] input_623;
    input [4:0] input_624;
    input [4:0] input_625;
    input [4:0] input_626;
    input [4:0] input_627;
    input [4:0] input_628;
    input [4:0] input_629;
    input [4:0] input_630;
    input [4:0] input_631;
    input [4:0] input_632;
    input [4:0] input_633;
    input [4:0] input_634;
    input [4:0] input_635;
    input [4:0] input_636;
    input [4:0] input_637;
    input [4:0] input_638;
    input [4:0] input_639;
    input [4:0] input_640;
    input [4:0] input_641;
    input [4:0] input_642;
    input [4:0] input_643;
    input [4:0] input_644;
    input [4:0] input_645;
    input [4:0] input_646;
    input [4:0] input_647;
    input [4:0] input_648;
    input [4:0] input_649;
    input [4:0] input_650;
    input [4:0] input_651;
    input [4:0] input_652;
    input [4:0] input_653;
    input [4:0] input_654;
    input [4:0] input_655;
    input [4:0] input_656;
    input [4:0] input_657;
    input [4:0] input_658;
    input [4:0] input_659;
    input [4:0] input_660;
    input [4:0] input_661;
    input [4:0] input_662;
    input [4:0] input_663;
    input [4:0] input_664;
    input [4:0] input_665;
    input [4:0] input_666;
    input [4:0] input_667;
    input [4:0] input_668;
    input [4:0] input_669;
    input [4:0] input_670;
    input [4:0] input_671;
    input [4:0] input_672;
    input [4:0] input_673;
    input [4:0] input_674;
    input [4:0] input_675;
    input [4:0] input_676;
    input [4:0] input_677;
    input [4:0] input_678;
    input [4:0] input_679;
    input [4:0] input_680;
    input [4:0] input_681;
    input [4:0] input_682;
    input [4:0] input_683;
    input [4:0] input_684;
    input [4:0] input_685;
    input [4:0] input_686;
    input [4:0] input_687;
    input [4:0] input_688;
    input [4:0] input_689;
    input [4:0] input_690;
    input [4:0] input_691;
    input [4:0] input_692;
    input [4:0] input_693;
    input [4:0] input_694;
    input [4:0] input_695;
    input [4:0] input_696;
    input [4:0] input_697;
    input [4:0] input_698;
    input [4:0] input_699;
    input [4:0] input_700;
    input [4:0] input_701;
    input [4:0] input_702;
    input [4:0] input_703;
    input [4:0] input_704;
    input [4:0] input_705;
    input [4:0] input_706;
    input [4:0] input_707;
    input [4:0] input_708;
    input [4:0] input_709;
    input [4:0] input_710;
    input [4:0] input_711;
    input [4:0] input_712;
    input [4:0] input_713;
    input [4:0] input_714;
    input [4:0] input_715;
    input [4:0] input_716;
    input [4:0] input_717;
    input [4:0] input_718;
    input [4:0] input_719;
    input [4:0] input_720;
    input [4:0] input_721;
    input [4:0] input_722;
    input [4:0] input_723;
    input [4:0] input_724;
    input [4:0] input_725;
    input [4:0] input_726;
    input [4:0] input_727;
    input [4:0] input_728;
    input [4:0] input_729;
    input [4:0] input_730;
    input [4:0] input_731;
    input [4:0] input_732;
    input [4:0] input_733;
    input [4:0] input_734;
    input [4:0] input_735;
    input [4:0] input_736;
    input [4:0] input_737;
    input [4:0] input_738;
    input [4:0] input_739;
    input [4:0] input_740;
    input [4:0] input_741;
    input [4:0] input_742;
    input [4:0] input_743;
    input [4:0] input_744;
    input [4:0] input_745;
    input [4:0] input_746;
    input [4:0] input_747;
    input [4:0] input_748;
    input [4:0] input_749;
    input [4:0] input_750;
    input [4:0] input_751;
    input [4:0] input_752;
    input [4:0] input_753;
    input [4:0] input_754;
    input [4:0] input_755;
    input [4:0] input_756;
    input [4:0] input_757;
    input [4:0] input_758;
    input [4:0] input_759;
    input [4:0] input_760;
    input [4:0] input_761;
    input [4:0] input_762;
    input [4:0] input_763;
    input [4:0] input_764;
    input [4:0] input_765;
    input [4:0] input_766;
    input [4:0] input_767;
    input [4:0] input_768;
    input [4:0] input_769;
    input [4:0] input_770;
    input [4:0] input_771;
    input [4:0] input_772;
    input [4:0] input_773;
    input [4:0] input_774;
    input [4:0] input_775;
    input [4:0] input_776;
    input [4:0] input_777;
    input [4:0] input_778;
    input [4:0] input_779;
    input [4:0] input_780;
    input [4:0] input_781;
    input [4:0] input_782;
    input [4:0] input_783;
    input [4:0] input_784;
    input [4:0] input_785;
    input [4:0] input_786;
    input [4:0] input_787;
    input [4:0] input_788;
    input [4:0] input_789;
    input [4:0] input_790;
    input [4:0] input_791;
    input [4:0] input_792;
    input [4:0] input_793;
    input [4:0] input_794;
    input [4:0] input_795;
    input [4:0] input_796;
    input [4:0] input_797;
    input [4:0] input_798;
    input [4:0] input_799;
    input [4:0] input_800;
    input [4:0] input_801;
    input [4:0] input_802;
    input [4:0] input_803;
    input [4:0] input_804;
    input [4:0] input_805;
    input [4:0] input_806;
    input [4:0] input_807;
    input [4:0] input_808;
    input [4:0] input_809;
    input [4:0] input_810;
    input [4:0] input_811;
    input [4:0] input_812;
    input [4:0] input_813;
    input [4:0] input_814;
    input [4:0] input_815;
    input [4:0] input_816;
    input [4:0] input_817;
    input [4:0] input_818;
    input [4:0] input_819;
    input [4:0] input_820;
    input [4:0] input_821;
    input [4:0] input_822;
    input [4:0] input_823;
    input [4:0] input_824;
    input [4:0] input_825;
    input [4:0] input_826;
    input [4:0] input_827;
    input [4:0] input_828;
    input [4:0] input_829;
    input [4:0] input_830;
    input [4:0] input_831;
    input [4:0] input_832;
    input [4:0] input_833;
    input [4:0] input_834;
    input [4:0] input_835;
    input [4:0] input_836;
    input [4:0] input_837;
    input [4:0] input_838;
    input [4:0] input_839;
    input [4:0] input_840;
    input [4:0] input_841;
    input [4:0] input_842;
    input [4:0] input_843;
    input [4:0] input_844;
    input [4:0] input_845;
    input [4:0] input_846;
    input [4:0] input_847;
    input [4:0] input_848;
    input [4:0] input_849;
    input [4:0] input_850;
    input [4:0] input_851;
    input [4:0] input_852;
    input [4:0] input_853;
    input [4:0] input_854;
    input [4:0] input_855;
    input [4:0] input_856;
    input [4:0] input_857;
    input [4:0] input_858;
    input [4:0] input_859;
    input [4:0] input_860;
    input [4:0] input_861;
    input [4:0] input_862;
    input [4:0] input_863;
    input [4:0] input_864;
    input [4:0] input_865;
    input [4:0] input_866;
    input [4:0] input_867;
    input [4:0] input_868;
    input [4:0] input_869;
    input [4:0] input_870;
    input [4:0] input_871;
    input [4:0] input_872;
    input [4:0] input_873;
    input [4:0] input_874;
    input [4:0] input_875;
    input [4:0] input_876;
    input [4:0] input_877;
    input [4:0] input_878;
    input [4:0] input_879;
    input [4:0] input_880;
    input [4:0] input_881;
    input [4:0] input_882;
    input [4:0] input_883;
    input [4:0] input_884;
    input [4:0] input_885;
    input [4:0] input_886;
    input [4:0] input_887;
    input [4:0] input_888;
    input [4:0] input_889;
    input [4:0] input_890;
    input [4:0] input_891;
    input [4:0] input_892;
    input [4:0] input_893;
    input [4:0] input_894;
    input [4:0] input_895;
    input [4:0] input_896;
    input [4:0] input_897;
    input [4:0] input_898;
    input [4:0] input_899;
    input [4:0] input_900;
    input [4:0] input_901;
    input [4:0] input_902;
    input [4:0] input_903;
    input [4:0] input_904;
    input [4:0] input_905;
    input [4:0] input_906;
    input [4:0] input_907;
    input [4:0] input_908;
    input [4:0] input_909;
    input [4:0] input_910;
    input [4:0] input_911;
    input [4:0] input_912;
    input [4:0] input_913;
    input [4:0] input_914;
    input [4:0] input_915;
    input [4:0] input_916;
    input [4:0] input_917;
    input [4:0] input_918;
    input [4:0] input_919;
    input [4:0] input_920;
    input [4:0] input_921;
    input [4:0] input_922;
    input [4:0] input_923;
    input [4:0] input_924;
    input [4:0] input_925;
    input [4:0] input_926;
    input [4:0] input_927;
    input [4:0] input_928;
    input [4:0] input_929;
    input [4:0] input_930;
    input [4:0] input_931;
    input [4:0] input_932;
    input [4:0] input_933;
    input [4:0] input_934;
    input [4:0] input_935;
    input [4:0] input_936;
    input [4:0] input_937;
    input [4:0] input_938;
    input [4:0] input_939;
    input [4:0] input_940;
    input [4:0] input_941;
    input [4:0] input_942;
    input [4:0] input_943;
    input [4:0] input_944;
    input [4:0] input_945;
    input [4:0] input_946;
    input [4:0] input_947;
    input [4:0] input_948;
    input [4:0] input_949;
    input [4:0] input_950;
    input [4:0] input_951;
    input [4:0] input_952;
    input [4:0] input_953;
    input [4:0] input_954;
    input [4:0] input_955;
    input [4:0] input_956;
    input [4:0] input_957;
    input [4:0] input_958;
    input [4:0] input_959;
    input [4:0] input_960;
    input [4:0] input_961;
    input [4:0] input_962;
    input [4:0] input_963;
    input [4:0] input_964;
    input [4:0] input_965;
    input [4:0] input_966;
    input [4:0] input_967;
    input [4:0] input_968;
    input [4:0] input_969;
    input [4:0] input_970;
    input [4:0] input_971;
    input [4:0] input_972;
    input [4:0] input_973;
    input [4:0] input_974;
    input [4:0] input_975;
    input [4:0] input_976;
    input [4:0] input_977;
    input [4:0] input_978;
    input [4:0] input_979;
    input [4:0] input_980;
    input [4:0] input_981;
    input [4:0] input_982;
    input [4:0] input_983;
    input [4:0] input_984;
    input [4:0] input_985;
    input [4:0] input_986;
    input [4:0] input_987;
    input [4:0] input_988;
    input [4:0] input_989;
    input [4:0] input_990;
    input [4:0] input_991;
    input [4:0] input_992;
    input [4:0] input_993;
    input [4:0] input_994;
    input [4:0] input_995;
    input [4:0] input_996;
    input [4:0] input_997;
    input [4:0] input_998;
    input [4:0] input_999;
    input [4:0] input_1000;
    input [4:0] input_1001;
    input [4:0] input_1002;
    input [4:0] input_1003;
    input [4:0] input_1004;
    input [4:0] input_1005;
    input [4:0] input_1006;
    input [4:0] input_1007;
    input [4:0] input_1008;
    input [4:0] input_1009;
    input [4:0] input_1010;
    input [4:0] input_1011;
    input [4:0] input_1012;
    input [4:0] input_1013;
    input [4:0] input_1014;
    input [4:0] input_1015;
    input [4:0] input_1016;
    input [4:0] input_1017;
    input [4:0] input_1018;
    input [4:0] input_1019;
    input [4:0] input_1020;
    input [4:0] input_1021;
    input [4:0] input_1022;
    input [4:0] input_1023;
    input [4:0] input_1024;
    input [4:0] input_1025;
    input [4:0] input_1026;
    input [4:0] input_1027;
    input [4:0] input_1028;
    input [4:0] input_1029;
    input [4:0] input_1030;
    input [4:0] input_1031;
    input [4:0] input_1032;
    input [4:0] input_1033;
    input [4:0] input_1034;
    input [4:0] input_1035;
    input [4:0] input_1036;
    input [4:0] input_1037;
    input [4:0] input_1038;
    input [4:0] input_1039;
    input [4:0] input_1040;
    input [4:0] input_1041;
    input [4:0] input_1042;
    input [4:0] input_1043;
    input [4:0] input_1044;
    input [4:0] input_1045;
    input [4:0] input_1046;
    input [4:0] input_1047;
    input [4:0] input_1048;
    input [4:0] input_1049;
    input [4:0] input_1050;
    input [4:0] input_1051;
    input [4:0] input_1052;
    input [4:0] input_1053;
    input [4:0] input_1054;
    input [4:0] input_1055;
    input [4:0] input_1056;
    input [4:0] input_1057;
    input [4:0] input_1058;
    input [4:0] input_1059;
    input [4:0] input_1060;
    input [4:0] input_1061;
    input [4:0] input_1062;
    input [4:0] input_1063;
    input [4:0] input_1064;
    input [4:0] input_1065;
    input [4:0] input_1066;
    input [4:0] input_1067;
    input [4:0] input_1068;
    input [4:0] input_1069;
    input [4:0] input_1070;
    input [4:0] input_1071;
    input [4:0] input_1072;
    input [4:0] input_1073;
    input [4:0] input_1074;
    input [4:0] input_1075;
    input [4:0] input_1076;
    input [4:0] input_1077;
    input [4:0] input_1078;
    input [4:0] input_1079;
    input [4:0] input_1080;
    input [4:0] input_1081;
    input [4:0] input_1082;
    input [4:0] input_1083;
    input [4:0] input_1084;
    input [4:0] input_1085;
    input [4:0] input_1086;
    input [4:0] input_1087;
    input [4:0] input_1088;
    input [4:0] input_1089;
    input [4:0] input_1090;
    input [4:0] input_1091;
    input [4:0] input_1092;
    input [4:0] input_1093;
    input [4:0] input_1094;
    input [4:0] input_1095;
    input [4:0] input_1096;
    input [4:0] input_1097;
    input [4:0] input_1098;
    input [4:0] input_1099;
    input [4:0] input_1100;
    input [4:0] input_1101;
    input [4:0] input_1102;
    input [4:0] input_1103;
    input [4:0] input_1104;
    input [4:0] input_1105;
    input [4:0] input_1106;
    input [4:0] input_1107;
    input [4:0] input_1108;
    input [4:0] input_1109;
    input [4:0] input_1110;
    input [4:0] input_1111;
    input [4:0] input_1112;
    input [4:0] input_1113;
    input [4:0] input_1114;
    input [4:0] input_1115;
    input [4:0] input_1116;
    input [4:0] input_1117;
    input [4:0] input_1118;
    input [4:0] input_1119;
    input [4:0] input_1120;
    input [4:0] input_1121;
    input [4:0] input_1122;
    input [4:0] input_1123;
    input [4:0] input_1124;
    input [4:0] input_1125;
    input [4:0] input_1126;
    input [4:0] input_1127;
    input [4:0] input_1128;
    input [4:0] input_1129;
    input [4:0] input_1130;
    input [4:0] input_1131;
    input [4:0] input_1132;
    input [4:0] input_1133;
    input [4:0] input_1134;
    input [4:0] input_1135;
    input [4:0] input_1136;
    input [4:0] input_1137;
    input [4:0] input_1138;
    input [4:0] input_1139;
    input [4:0] input_1140;
    input [4:0] input_1141;
    input [4:0] input_1142;
    input [4:0] input_1143;
    input [4:0] input_1144;
    input [4:0] input_1145;
    input [4:0] input_1146;
    input [4:0] input_1147;
    input [4:0] input_1148;
    input [4:0] input_1149;
    input [4:0] input_1150;
    input [4:0] input_1151;
    input [4:0] input_1152;
    input [4:0] input_1153;
    input [4:0] input_1154;
    input [4:0] input_1155;
    input [4:0] input_1156;
    input [4:0] input_1157;
    input [4:0] input_1158;
    input [4:0] input_1159;
    input [4:0] input_1160;
    input [4:0] input_1161;
    input [4:0] input_1162;
    input [4:0] input_1163;
    input [4:0] input_1164;
    input [4:0] input_1165;
    input [4:0] input_1166;
    input [4:0] input_1167;
    input [4:0] input_1168;
    input [4:0] input_1169;
    input [4:0] input_1170;
    input [4:0] input_1171;
    input [4:0] input_1172;
    input [4:0] input_1173;
    input [4:0] input_1174;
    input [4:0] input_1175;
    input [4:0] input_1176;
    input [4:0] input_1177;
    input [4:0] input_1178;
    input [4:0] input_1179;
    input [4:0] input_1180;
    input [4:0] input_1181;
    input [4:0] input_1182;
    input [4:0] input_1183;
    input [4:0] input_1184;
    input [4:0] input_1185;
    input [4:0] input_1186;
    input [4:0] input_1187;
    input [4:0] input_1188;
    input [4:0] input_1189;
    input [4:0] input_1190;
    input [4:0] input_1191;
    input [4:0] input_1192;
    input [4:0] input_1193;
    input [4:0] input_1194;
    input [4:0] input_1195;
    input [4:0] input_1196;
    input [4:0] input_1197;
    input [4:0] input_1198;
    input [4:0] input_1199;
    input [4:0] input_1200;
    input [4:0] input_1201;
    input [4:0] input_1202;
    input [4:0] input_1203;
    input [4:0] input_1204;
    input [4:0] input_1205;
    input [4:0] input_1206;
    input [4:0] input_1207;
    input [4:0] input_1208;
    input [4:0] input_1209;
    input [4:0] input_1210;
    input [4:0] input_1211;
    input [4:0] input_1212;
    input [4:0] input_1213;
    input [4:0] input_1214;
    input [4:0] input_1215;
    input [4:0] input_1216;
    input [4:0] input_1217;
    input [4:0] input_1218;
    input [4:0] input_1219;
    input [4:0] input_1220;
    input [4:0] input_1221;
    input [4:0] input_1222;
    input [4:0] input_1223;
    input [4:0] input_1224;
    input [4:0] input_1225;
    input [4:0] input_1226;
    input [4:0] input_1227;
    input [4:0] input_1228;
    input [4:0] input_1229;
    input [4:0] input_1230;
    input [4:0] input_1231;
    input [4:0] input_1232;
    input [4:0] input_1233;
    input [4:0] input_1234;
    input [4:0] input_1235;
    input [4:0] input_1236;
    input [4:0] input_1237;
    input [4:0] input_1238;
    input [4:0] input_1239;
    input [4:0] input_1240;
    input [4:0] input_1241;
    input [4:0] input_1242;
    input [4:0] input_1243;
    input [4:0] input_1244;
    input [4:0] input_1245;
    input [4:0] input_1246;
    input [4:0] input_1247;
    input [4:0] input_1248;
    input [4:0] input_1249;
    input [4:0] input_1250;
    input [4:0] input_1251;
    input [4:0] input_1252;
    input [4:0] input_1253;
    input [4:0] input_1254;
    input [4:0] input_1255;
    input [4:0] input_1256;
    input [4:0] input_1257;
    input [4:0] input_1258;
    input [4:0] input_1259;
    input [4:0] input_1260;
    input [4:0] input_1261;
    input [4:0] input_1262;
    input [4:0] input_1263;
    input [4:0] input_1264;
    input [4:0] input_1265;
    input [4:0] input_1266;
    input [4:0] input_1267;
    input [4:0] input_1268;
    input [4:0] input_1269;
    input [4:0] input_1270;
    input [4:0] input_1271;
    input [4:0] input_1272;
    input [4:0] input_1273;
    input [4:0] input_1274;
    input [4:0] input_1275;
    input [4:0] input_1276;
    input [4:0] input_1277;
    input [4:0] input_1278;
    input [4:0] input_1279;
    input [4:0] input_1280;
    input [4:0] input_1281;
    input [4:0] input_1282;
    input [4:0] input_1283;
    input [4:0] input_1284;
    input [4:0] input_1285;
    input [4:0] input_1286;
    input [4:0] input_1287;
    input [4:0] input_1288;
    input [4:0] input_1289;
    input [4:0] input_1290;
    input [4:0] input_1291;
    input [4:0] input_1292;
    input [4:0] input_1293;
    input [4:0] input_1294;
    input [4:0] input_1295;
    input [4:0] input_1296;
    input [4:0] input_1297;
    input [4:0] input_1298;
    input [4:0] input_1299;
    input [4:0] input_1300;
    input [4:0] input_1301;
    input [4:0] input_1302;
    input [4:0] input_1303;
    input [4:0] input_1304;
    input [4:0] input_1305;
    input [4:0] input_1306;
    input [4:0] input_1307;
    input [4:0] input_1308;
    input [4:0] input_1309;
    input [4:0] input_1310;
    input [4:0] input_1311;
    input [4:0] input_1312;
    input [4:0] input_1313;
    input [4:0] input_1314;
    input [4:0] input_1315;
    input [4:0] input_1316;
    input [4:0] input_1317;
    input [4:0] input_1318;
    input [4:0] input_1319;
    input [4:0] input_1320;
    input [4:0] input_1321;
    input [4:0] input_1322;
    input [4:0] input_1323;
    input [4:0] input_1324;
    input [4:0] input_1325;
    input [4:0] input_1326;
    input [4:0] input_1327;
    input [4:0] input_1328;
    input [4:0] input_1329;
    input [4:0] input_1330;
    input [4:0] input_1331;
    input [4:0] input_1332;
    input [4:0] input_1333;
    input [4:0] input_1334;
    input [4:0] input_1335;
    input [4:0] input_1336;
    input [4:0] input_1337;
    input [4:0] input_1338;
    input [4:0] input_1339;
    input [4:0] input_1340;
    input [4:0] input_1341;
    input [4:0] input_1342;
    input [4:0] input_1343;
    input [4:0] input_1344;
    input [4:0] input_1345;
    input [4:0] input_1346;
    input [4:0] input_1347;
    input [4:0] input_1348;
    input [4:0] input_1349;
    input [4:0] input_1350;
    input [4:0] input_1351;
    input [4:0] input_1352;
    input [4:0] input_1353;
    input [4:0] input_1354;
    input [4:0] input_1355;
    input [4:0] input_1356;
    input [4:0] input_1357;
    input [4:0] input_1358;
    input [4:0] input_1359;
    input [4:0] input_1360;
    input [4:0] input_1361;
    input [4:0] input_1362;
    input [4:0] input_1363;
    input [4:0] input_1364;
    input [4:0] input_1365;
    input [4:0] input_1366;
    input [4:0] input_1367;
    input [4:0] input_1368;
    input [4:0] input_1369;
    input [4:0] input_1370;
    input [4:0] input_1371;
    input [4:0] input_1372;
    input [4:0] input_1373;
    input [4:0] input_1374;
    input [4:0] input_1375;
    input [4:0] input_1376;
    input [4:0] input_1377;
    input [4:0] input_1378;
    input [4:0] input_1379;
    input [4:0] input_1380;
    input [4:0] input_1381;
    input [4:0] input_1382;
    input [4:0] input_1383;
    input [4:0] input_1384;
    input [4:0] input_1385;
    input [4:0] input_1386;
    input [4:0] input_1387;
    input [4:0] input_1388;
    input [4:0] input_1389;
    input [4:0] input_1390;
    input [4:0] input_1391;
    input [4:0] input_1392;
    input [4:0] input_1393;
    input [4:0] input_1394;
    input [4:0] input_1395;
    input [4:0] input_1396;
    input [4:0] input_1397;
    input [4:0] input_1398;
    input [4:0] input_1399;
    input [4:0] input_1400;
    input [4:0] input_1401;
    input [4:0] input_1402;
    input [4:0] input_1403;
    input [4:0] input_1404;
    input [4:0] input_1405;
    input [4:0] input_1406;
    input [4:0] input_1407;
    input [4:0] input_1408;
    input [4:0] input_1409;
    input [4:0] input_1410;
    input [4:0] input_1411;
    input [4:0] input_1412;
    input [4:0] input_1413;
    input [4:0] input_1414;
    input [4:0] input_1415;
    input [4:0] input_1416;
    input [4:0] input_1417;
    input [4:0] input_1418;
    input [4:0] input_1419;
    input [4:0] input_1420;
    input [4:0] input_1421;
    input [4:0] input_1422;
    input [4:0] input_1423;
    input [4:0] input_1424;
    input [4:0] input_1425;
    input [4:0] input_1426;
    input [4:0] input_1427;
    input [4:0] input_1428;
    input [4:0] input_1429;
    input [4:0] input_1430;
    input [4:0] input_1431;
    input [4:0] input_1432;
    input [4:0] input_1433;
    input [4:0] input_1434;
    input [4:0] input_1435;
    input [4:0] input_1436;
    input [4:0] input_1437;
    input [4:0] input_1438;
    input [4:0] input_1439;
    input [4:0] input_1440;
    input [4:0] input_1441;
    input [4:0] input_1442;
    input [4:0] input_1443;
    input [4:0] input_1444;
    input [4:0] input_1445;
    input [4:0] input_1446;
    input [4:0] input_1447;
    input [4:0] input_1448;
    input [4:0] input_1449;
    input [4:0] input_1450;
    input [4:0] input_1451;
    input [4:0] input_1452;
    input [4:0] input_1453;
    input [4:0] input_1454;
    input [4:0] input_1455;
    input [4:0] input_1456;
    input [4:0] input_1457;
    input [4:0] input_1458;
    input [4:0] input_1459;
    input [4:0] input_1460;
    input [4:0] input_1461;
    input [4:0] input_1462;
    input [4:0] input_1463;
    input [4:0] input_1464;
    input [4:0] input_1465;
    input [4:0] input_1466;
    input [4:0] input_1467;
    input [4:0] input_1468;
    input [4:0] input_1469;
    input [4:0] input_1470;
    input [4:0] input_1471;
    input [4:0] input_1472;
    input [4:0] input_1473;
    input [4:0] input_1474;
    input [4:0] input_1475;
    input [4:0] input_1476;
    input [4:0] input_1477;
    input [4:0] input_1478;
    input [4:0] input_1479;
    input [4:0] input_1480;
    input [4:0] input_1481;
    input [4:0] input_1482;
    input [4:0] input_1483;
    input [4:0] input_1484;
    input [4:0] input_1485;
    input [4:0] input_1486;
    input [4:0] input_1487;
    input [4:0] input_1488;
    input [4:0] input_1489;
    input [4:0] input_1490;
    input [4:0] input_1491;
    input [4:0] input_1492;
    input [4:0] input_1493;
    input [4:0] input_1494;
    input [4:0] input_1495;
    input [4:0] input_1496;
    input [4:0] input_1497;
    input [4:0] input_1498;
    input [4:0] input_1499;
    input [4:0] input_1500;
    input [4:0] input_1501;
    input [4:0] input_1502;
    input [4:0] input_1503;
    input [4:0] input_1504;
    input [4:0] input_1505;
    input [4:0] input_1506;
    input [4:0] input_1507;
    input [4:0] input_1508;
    input [4:0] input_1509;
    input [4:0] input_1510;
    input [4:0] input_1511;
    input [4:0] input_1512;
    input [4:0] input_1513;
    input [4:0] input_1514;
    input [4:0] input_1515;
    input [4:0] input_1516;
    input [4:0] input_1517;
    input [4:0] input_1518;
    input [4:0] input_1519;
    input [4:0] input_1520;
    input [4:0] input_1521;
    input [4:0] input_1522;
    input [4:0] input_1523;
    input [4:0] input_1524;
    input [4:0] input_1525;
    input [4:0] input_1526;
    input [4:0] input_1527;
    input [4:0] input_1528;
    input [4:0] input_1529;
    input [4:0] input_1530;
    input [4:0] input_1531;
    input [4:0] input_1532;
    input [4:0] input_1533;
    input [4:0] input_1534;
    input [4:0] input_1535;
    input [4:0] input_1536;
    input [4:0] input_1537;
    input [4:0] input_1538;
    input [4:0] input_1539;
    input [4:0] input_1540;
    input [4:0] input_1541;
    input [4:0] input_1542;
    input [4:0] input_1543;
    input [4:0] input_1544;
    input [4:0] input_1545;
    input [4:0] input_1546;
    input [4:0] input_1547;
    input [4:0] input_1548;
    input [4:0] input_1549;
    input [4:0] input_1550;
    input [4:0] input_1551;
    input [4:0] input_1552;
    input [4:0] input_1553;
    input [4:0] input_1554;
    input [4:0] input_1555;
    input [4:0] input_1556;
    input [4:0] input_1557;
    input [4:0] input_1558;
    input [4:0] input_1559;
    input [4:0] input_1560;
    input [4:0] input_1561;
    input [4:0] input_1562;
    input [4:0] input_1563;
    input [4:0] input_1564;
    input [4:0] input_1565;
    input [4:0] input_1566;
    input [4:0] input_1567;
    input [4:0] input_1568;
    input [4:0] input_1569;
    input [4:0] input_1570;
    input [4:0] input_1571;
    input [4:0] input_1572;
    input [4:0] input_1573;
    input [4:0] input_1574;
    input [4:0] input_1575;
    input [4:0] input_1576;
    input [4:0] input_1577;
    input [4:0] input_1578;
    input [4:0] input_1579;
    input [4:0] input_1580;
    input [4:0] input_1581;
    input [4:0] input_1582;
    input [4:0] input_1583;
    input [4:0] input_1584;
    input [4:0] input_1585;
    input [4:0] input_1586;
    input [4:0] input_1587;
    input [4:0] input_1588;
    input [4:0] input_1589;
    input [4:0] input_1590;
    input [4:0] input_1591;
    input [4:0] input_1592;
    input [4:0] input_1593;
    input [4:0] input_1594;
    input [4:0] input_1595;
    input [4:0] input_1596;
    input [4:0] input_1597;
    input [4:0] input_1598;
    input [4:0] input_1599;
    input [4:0] input_1600;
    input [4:0] input_1601;
    input [4:0] input_1602;
    input [4:0] input_1603;
    input [4:0] input_1604;
    input [4:0] input_1605;
    input [4:0] input_1606;
    input [4:0] input_1607;
    input [4:0] input_1608;
    input [4:0] input_1609;
    input [4:0] input_1610;
    input [4:0] input_1611;
    input [4:0] input_1612;
    input [4:0] input_1613;
    input [4:0] input_1614;
    input [4:0] input_1615;
    input [4:0] input_1616;
    input [4:0] input_1617;
    input [4:0] input_1618;
    input [4:0] input_1619;
    input [4:0] input_1620;
    input [4:0] input_1621;
    input [4:0] input_1622;
    input [4:0] input_1623;
    input [4:0] input_1624;
    input [4:0] input_1625;
    input [4:0] input_1626;
    input [4:0] input_1627;
    input [4:0] input_1628;
    input [4:0] input_1629;
    input [4:0] input_1630;
    input [4:0] input_1631;
    input [4:0] input_1632;
    input [4:0] input_1633;
    input [4:0] input_1634;
    input [4:0] input_1635;
    input [4:0] input_1636;
    input [4:0] input_1637;
    input [4:0] input_1638;
    input [4:0] input_1639;
    input [4:0] input_1640;
    input [4:0] input_1641;
    input [4:0] input_1642;
    input [4:0] input_1643;
    input [4:0] input_1644;
    input [4:0] input_1645;
    input [4:0] input_1646;
    input [4:0] input_1647;
    input [4:0] input_1648;
    input [4:0] input_1649;
    input [4:0] input_1650;
    input [4:0] input_1651;
    input [4:0] input_1652;
    input [4:0] input_1653;
    input [4:0] input_1654;
    input [4:0] input_1655;
    input [4:0] input_1656;
    input [4:0] input_1657;
    input [4:0] input_1658;
    input [4:0] input_1659;
    input [4:0] input_1660;
    input [4:0] input_1661;
    input [4:0] input_1662;
    input [4:0] input_1663;
    input [4:0] input_1664;
    input [4:0] input_1665;
    input [4:0] input_1666;
    input [4:0] input_1667;
    input [4:0] input_1668;
    input [4:0] input_1669;
    input [4:0] input_1670;
    input [4:0] input_1671;
    input [4:0] input_1672;
    input [4:0] input_1673;
    input [4:0] input_1674;
    input [4:0] input_1675;
    input [4:0] input_1676;
    input [4:0] input_1677;
    input [4:0] input_1678;
    input [4:0] input_1679;
    input [4:0] input_1680;
    input [4:0] input_1681;
    input [4:0] input_1682;
    input [4:0] input_1683;
    input [4:0] input_1684;
    input [4:0] input_1685;
    input [4:0] input_1686;
    input [4:0] input_1687;
    input [4:0] input_1688;
    input [4:0] input_1689;
    input [4:0] input_1690;
    input [4:0] input_1691;
    input [4:0] input_1692;
    input [4:0] input_1693;
    input [4:0] input_1694;
    input [4:0] input_1695;
    input [4:0] input_1696;
    input [4:0] input_1697;
    input [4:0] input_1698;
    input [4:0] input_1699;
    input [4:0] input_1700;
    input [4:0] input_1701;
    input [4:0] input_1702;
    input [4:0] input_1703;
    input [4:0] input_1704;
    input [4:0] input_1705;
    input [4:0] input_1706;
    input [4:0] input_1707;
    input [4:0] input_1708;
    input [4:0] input_1709;
    input [4:0] input_1710;
    input [4:0] input_1711;
    input [4:0] input_1712;
    input [4:0] input_1713;
    input [4:0] input_1714;
    input [4:0] input_1715;
    input [4:0] input_1716;
    input [4:0] input_1717;
    input [4:0] input_1718;
    input [4:0] input_1719;
    input [4:0] input_1720;
    input [4:0] input_1721;
    input [4:0] input_1722;
    input [4:0] input_1723;
    input [4:0] input_1724;
    input [4:0] input_1725;
    input [4:0] input_1726;
    input [4:0] input_1727;
    input [4:0] input_1728;
    input [4:0] input_1729;
    input [4:0] input_1730;
    input [4:0] input_1731;
    input [4:0] input_1732;
    input [4:0] input_1733;
    input [4:0] input_1734;
    input [4:0] input_1735;
    input [4:0] input_1736;
    input [4:0] input_1737;
    input [4:0] input_1738;
    input [4:0] input_1739;
    input [4:0] input_1740;
    input [4:0] input_1741;
    input [4:0] input_1742;
    input [4:0] input_1743;
    input [4:0] input_1744;
    input [4:0] input_1745;
    input [4:0] input_1746;
    input [4:0] input_1747;
    input [4:0] input_1748;
    input [4:0] input_1749;
    input [4:0] input_1750;
    input [4:0] input_1751;
    input [4:0] input_1752;
    input [4:0] input_1753;
    input [4:0] input_1754;
    input [4:0] input_1755;
    input [4:0] input_1756;
    input [4:0] input_1757;
    input [4:0] input_1758;
    input [4:0] input_1759;
    input [4:0] input_1760;
    input [4:0] input_1761;
    input [4:0] input_1762;
    input [4:0] input_1763;
    input [4:0] input_1764;
    input [4:0] input_1765;
    input [4:0] input_1766;
    input [4:0] input_1767;
    input [4:0] input_1768;
    input [4:0] input_1769;
    input [4:0] input_1770;
    input [4:0] input_1771;
    input [4:0] input_1772;
    input [4:0] input_1773;
    input [4:0] input_1774;
    input [4:0] input_1775;
    input [4:0] input_1776;
    input [4:0] input_1777;
    input [4:0] input_1778;
    input [4:0] input_1779;
    input [4:0] input_1780;
    input [4:0] input_1781;
    input [4:0] input_1782;
    input [4:0] input_1783;
    input [4:0] input_1784;
    input [4:0] input_1785;
    input [4:0] input_1786;
    input [4:0] input_1787;
    input [4:0] input_1788;
    input [4:0] input_1789;
    input [4:0] input_1790;
    input [4:0] input_1791;
    input [4:0] input_1792;
    input [4:0] input_1793;
    input [4:0] input_1794;
    input [4:0] input_1795;
    input [4:0] input_1796;
    input [4:0] input_1797;
    input [4:0] input_1798;
    input [4:0] input_1799;
    input [4:0] input_1800;
    input [4:0] input_1801;
    input [4:0] input_1802;
    input [4:0] input_1803;
    input [4:0] input_1804;
    input [4:0] input_1805;
    input [4:0] input_1806;
    input [4:0] input_1807;
    input [4:0] input_1808;
    input [4:0] input_1809;
    input [4:0] input_1810;
    input [4:0] input_1811;
    input [4:0] input_1812;
    input [4:0] input_1813;
    input [4:0] input_1814;
    input [4:0] input_1815;
    input [4:0] input_1816;
    input [4:0] input_1817;
    input [4:0] input_1818;
    input [4:0] input_1819;
    input [4:0] input_1820;
    input [4:0] input_1821;
    input [4:0] input_1822;
    input [4:0] input_1823;
    input [4:0] input_1824;
    input [4:0] input_1825;
    input [4:0] input_1826;
    input [4:0] input_1827;
    input [4:0] input_1828;
    input [4:0] input_1829;
    input [4:0] input_1830;
    input [4:0] input_1831;
    input [4:0] input_1832;
    input [4:0] input_1833;
    input [4:0] input_1834;
    input [4:0] input_1835;
    input [4:0] input_1836;
    input [4:0] input_1837;
    input [4:0] input_1838;
    input [4:0] input_1839;
    input [4:0] input_1840;
    input [4:0] input_1841;
    input [4:0] input_1842;
    input [4:0] input_1843;
    input [4:0] input_1844;
    input [4:0] input_1845;
    input [4:0] input_1846;
    input [4:0] input_1847;
    input [4:0] input_1848;
    input [4:0] input_1849;
    input [4:0] input_1850;
    input [4:0] input_1851;
    input [4:0] input_1852;
    input [4:0] input_1853;
    input [4:0] input_1854;
    input [4:0] input_1855;
    input [4:0] input_1856;
    input [4:0] input_1857;
    input [4:0] input_1858;
    input [4:0] input_1859;
    input [4:0] input_1860;
    input [4:0] input_1861;
    input [4:0] input_1862;
    input [4:0] input_1863;
    input [4:0] input_1864;
    input [4:0] input_1865;
    input [4:0] input_1866;
    input [4:0] input_1867;
    input [4:0] input_1868;
    input [4:0] input_1869;
    input [4:0] input_1870;
    input [4:0] input_1871;
    input [4:0] input_1872;
    input [4:0] input_1873;
    input [4:0] input_1874;
    input [4:0] input_1875;
    input [4:0] input_1876;
    input [4:0] input_1877;
    input [4:0] input_1878;
    input [4:0] input_1879;
    input [4:0] input_1880;
    input [4:0] input_1881;
    input [4:0] input_1882;
    input [4:0] input_1883;
    input [4:0] input_1884;
    input [4:0] input_1885;
    input [4:0] input_1886;
    input [4:0] input_1887;
    input [4:0] input_1888;
    input [4:0] input_1889;
    input [4:0] input_1890;
    input [4:0] input_1891;
    input [4:0] input_1892;
    input [4:0] input_1893;
    input [4:0] input_1894;
    input [4:0] input_1895;
    input [4:0] input_1896;
    input [4:0] input_1897;
    input [4:0] input_1898;
    input [4:0] input_1899;
    input [4:0] input_1900;
    input [4:0] input_1901;
    input [4:0] input_1902;
    input [4:0] input_1903;
    input [4:0] input_1904;
    input [4:0] input_1905;
    input [4:0] input_1906;
    input [4:0] input_1907;
    input [4:0] input_1908;
    input [4:0] input_1909;
    input [4:0] input_1910;
    input [4:0] input_1911;
    input [4:0] input_1912;
    input [4:0] input_1913;
    input [4:0] input_1914;
    input [4:0] input_1915;
    input [4:0] input_1916;
    input [4:0] input_1917;
    input [4:0] input_1918;
    input [4:0] input_1919;
    input [4:0] input_1920;
    input [4:0] input_1921;
    input [4:0] input_1922;
    input [4:0] input_1923;
    input [4:0] input_1924;
    input [4:0] input_1925;
    input [4:0] input_1926;
    input [4:0] input_1927;
    input [4:0] input_1928;
    input [4:0] input_1929;
    input [4:0] input_1930;
    input [4:0] input_1931;
    input [4:0] input_1932;
    input [4:0] input_1933;
    input [4:0] input_1934;
    input [4:0] input_1935;
    input [4:0] input_1936;
    input [4:0] input_1937;
    input [4:0] input_1938;
    input [4:0] input_1939;
    input [4:0] input_1940;
    input [4:0] input_1941;
    input [4:0] input_1942;
    input [4:0] input_1943;
    input [4:0] input_1944;
    input [4:0] input_1945;
    input [4:0] input_1946;
    input [4:0] input_1947;
    input [4:0] input_1948;
    input [4:0] input_1949;
    input [4:0] input_1950;
    input [4:0] input_1951;
    input [4:0] input_1952;
    input [4:0] input_1953;
    input [4:0] input_1954;
    input [4:0] input_1955;
    input [4:0] input_1956;
    input [4:0] input_1957;
    input [4:0] input_1958;
    input [4:0] input_1959;
    input [4:0] input_1960;
    input [4:0] input_1961;
    input [4:0] input_1962;
    input [4:0] input_1963;
    input [4:0] input_1964;
    input [4:0] input_1965;
    input [4:0] input_1966;
    input [4:0] input_1967;
    input [4:0] input_1968;
    input [4:0] input_1969;
    input [4:0] input_1970;
    input [4:0] input_1971;
    input [4:0] input_1972;
    input [4:0] input_1973;
    input [4:0] input_1974;
    input [4:0] input_1975;
    input [4:0] input_1976;
    input [4:0] input_1977;
    input [4:0] input_1978;
    input [4:0] input_1979;
    input [4:0] input_1980;
    input [4:0] input_1981;
    input [4:0] input_1982;
    input [4:0] input_1983;
    input [4:0] input_1984;
    input [4:0] input_1985;
    input [4:0] input_1986;
    input [4:0] input_1987;
    input [4:0] input_1988;
    input [4:0] input_1989;
    input [4:0] input_1990;
    input [4:0] input_1991;
    input [4:0] input_1992;
    input [4:0] input_1993;
    input [4:0] input_1994;
    input [4:0] input_1995;
    input [4:0] input_1996;
    input [4:0] input_1997;
    input [4:0] input_1998;
    input [4:0] input_1999;
    input [4:0] input_2000;
    input [4:0] input_2001;
    input [4:0] input_2002;
    input [4:0] input_2003;
    input [4:0] input_2004;
    input [4:0] input_2005;
    input [4:0] input_2006;
    input [4:0] input_2007;
    input [4:0] input_2008;
    input [4:0] input_2009;
    input [4:0] input_2010;
    input [4:0] input_2011;
    input [4:0] input_2012;
    input [4:0] input_2013;
    input [4:0] input_2014;
    input [4:0] input_2015;
    input [4:0] input_2016;
    input [4:0] input_2017;
    input [4:0] input_2018;
    input [4:0] input_2019;
    input [4:0] input_2020;
    input [4:0] input_2021;
    input [4:0] input_2022;
    input [4:0] input_2023;
    input [4:0] input_2024;
    input [4:0] input_2025;
    input [4:0] input_2026;
    input [4:0] input_2027;
    input [4:0] input_2028;
    input [4:0] input_2029;
    input [4:0] input_2030;
    input [4:0] input_2031;
    input [4:0] input_2032;
    input [4:0] input_2033;
    input [4:0] input_2034;
    input [4:0] input_2035;
    input [4:0] input_2036;
    input [4:0] input_2037;
    input [4:0] input_2038;
    input [4:0] input_2039;
    input [4:0] input_2040;
    input [4:0] input_2041;
    input [4:0] input_2042;
    input [4:0] input_2043;
    input [4:0] input_2044;
    input [4:0] input_2045;
    input [4:0] input_2046;
    input [4:0] input_2047;
    input [10:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      11'b00000000000 : begin
        result = input_0;
      end
      11'b00000000001 : begin
        result = input_1;
      end
      11'b00000000010 : begin
        result = input_2;
      end
      11'b00000000011 : begin
        result = input_3;
      end
      11'b00000000100 : begin
        result = input_4;
      end
      11'b00000000101 : begin
        result = input_5;
      end
      11'b00000000110 : begin
        result = input_6;
      end
      11'b00000000111 : begin
        result = input_7;
      end
      11'b00000001000 : begin
        result = input_8;
      end
      11'b00000001001 : begin
        result = input_9;
      end
      11'b00000001010 : begin
        result = input_10;
      end
      11'b00000001011 : begin
        result = input_11;
      end
      11'b00000001100 : begin
        result = input_12;
      end
      11'b00000001101 : begin
        result = input_13;
      end
      11'b00000001110 : begin
        result = input_14;
      end
      11'b00000001111 : begin
        result = input_15;
      end
      11'b00000010000 : begin
        result = input_16;
      end
      11'b00000010001 : begin
        result = input_17;
      end
      11'b00000010010 : begin
        result = input_18;
      end
      11'b00000010011 : begin
        result = input_19;
      end
      11'b00000010100 : begin
        result = input_20;
      end
      11'b00000010101 : begin
        result = input_21;
      end
      11'b00000010110 : begin
        result = input_22;
      end
      11'b00000010111 : begin
        result = input_23;
      end
      11'b00000011000 : begin
        result = input_24;
      end
      11'b00000011001 : begin
        result = input_25;
      end
      11'b00000011010 : begin
        result = input_26;
      end
      11'b00000011011 : begin
        result = input_27;
      end
      11'b00000011100 : begin
        result = input_28;
      end
      11'b00000011101 : begin
        result = input_29;
      end
      11'b00000011110 : begin
        result = input_30;
      end
      11'b00000011111 : begin
        result = input_31;
      end
      11'b00000100000 : begin
        result = input_32;
      end
      11'b00000100001 : begin
        result = input_33;
      end
      11'b00000100010 : begin
        result = input_34;
      end
      11'b00000100011 : begin
        result = input_35;
      end
      11'b00000100100 : begin
        result = input_36;
      end
      11'b00000100101 : begin
        result = input_37;
      end
      11'b00000100110 : begin
        result = input_38;
      end
      11'b00000100111 : begin
        result = input_39;
      end
      11'b00000101000 : begin
        result = input_40;
      end
      11'b00000101001 : begin
        result = input_41;
      end
      11'b00000101010 : begin
        result = input_42;
      end
      11'b00000101011 : begin
        result = input_43;
      end
      11'b00000101100 : begin
        result = input_44;
      end
      11'b00000101101 : begin
        result = input_45;
      end
      11'b00000101110 : begin
        result = input_46;
      end
      11'b00000101111 : begin
        result = input_47;
      end
      11'b00000110000 : begin
        result = input_48;
      end
      11'b00000110001 : begin
        result = input_49;
      end
      11'b00000110010 : begin
        result = input_50;
      end
      11'b00000110011 : begin
        result = input_51;
      end
      11'b00000110100 : begin
        result = input_52;
      end
      11'b00000110101 : begin
        result = input_53;
      end
      11'b00000110110 : begin
        result = input_54;
      end
      11'b00000110111 : begin
        result = input_55;
      end
      11'b00000111000 : begin
        result = input_56;
      end
      11'b00000111001 : begin
        result = input_57;
      end
      11'b00000111010 : begin
        result = input_58;
      end
      11'b00000111011 : begin
        result = input_59;
      end
      11'b00000111100 : begin
        result = input_60;
      end
      11'b00000111101 : begin
        result = input_61;
      end
      11'b00000111110 : begin
        result = input_62;
      end
      11'b00000111111 : begin
        result = input_63;
      end
      11'b00001000000 : begin
        result = input_64;
      end
      11'b00001000001 : begin
        result = input_65;
      end
      11'b00001000010 : begin
        result = input_66;
      end
      11'b00001000011 : begin
        result = input_67;
      end
      11'b00001000100 : begin
        result = input_68;
      end
      11'b00001000101 : begin
        result = input_69;
      end
      11'b00001000110 : begin
        result = input_70;
      end
      11'b00001000111 : begin
        result = input_71;
      end
      11'b00001001000 : begin
        result = input_72;
      end
      11'b00001001001 : begin
        result = input_73;
      end
      11'b00001001010 : begin
        result = input_74;
      end
      11'b00001001011 : begin
        result = input_75;
      end
      11'b00001001100 : begin
        result = input_76;
      end
      11'b00001001101 : begin
        result = input_77;
      end
      11'b00001001110 : begin
        result = input_78;
      end
      11'b00001001111 : begin
        result = input_79;
      end
      11'b00001010000 : begin
        result = input_80;
      end
      11'b00001010001 : begin
        result = input_81;
      end
      11'b00001010010 : begin
        result = input_82;
      end
      11'b00001010011 : begin
        result = input_83;
      end
      11'b00001010100 : begin
        result = input_84;
      end
      11'b00001010101 : begin
        result = input_85;
      end
      11'b00001010110 : begin
        result = input_86;
      end
      11'b00001010111 : begin
        result = input_87;
      end
      11'b00001011000 : begin
        result = input_88;
      end
      11'b00001011001 : begin
        result = input_89;
      end
      11'b00001011010 : begin
        result = input_90;
      end
      11'b00001011011 : begin
        result = input_91;
      end
      11'b00001011100 : begin
        result = input_92;
      end
      11'b00001011101 : begin
        result = input_93;
      end
      11'b00001011110 : begin
        result = input_94;
      end
      11'b00001011111 : begin
        result = input_95;
      end
      11'b00001100000 : begin
        result = input_96;
      end
      11'b00001100001 : begin
        result = input_97;
      end
      11'b00001100010 : begin
        result = input_98;
      end
      11'b00001100011 : begin
        result = input_99;
      end
      11'b00001100100 : begin
        result = input_100;
      end
      11'b00001100101 : begin
        result = input_101;
      end
      11'b00001100110 : begin
        result = input_102;
      end
      11'b00001100111 : begin
        result = input_103;
      end
      11'b00001101000 : begin
        result = input_104;
      end
      11'b00001101001 : begin
        result = input_105;
      end
      11'b00001101010 : begin
        result = input_106;
      end
      11'b00001101011 : begin
        result = input_107;
      end
      11'b00001101100 : begin
        result = input_108;
      end
      11'b00001101101 : begin
        result = input_109;
      end
      11'b00001101110 : begin
        result = input_110;
      end
      11'b00001101111 : begin
        result = input_111;
      end
      11'b00001110000 : begin
        result = input_112;
      end
      11'b00001110001 : begin
        result = input_113;
      end
      11'b00001110010 : begin
        result = input_114;
      end
      11'b00001110011 : begin
        result = input_115;
      end
      11'b00001110100 : begin
        result = input_116;
      end
      11'b00001110101 : begin
        result = input_117;
      end
      11'b00001110110 : begin
        result = input_118;
      end
      11'b00001110111 : begin
        result = input_119;
      end
      11'b00001111000 : begin
        result = input_120;
      end
      11'b00001111001 : begin
        result = input_121;
      end
      11'b00001111010 : begin
        result = input_122;
      end
      11'b00001111011 : begin
        result = input_123;
      end
      11'b00001111100 : begin
        result = input_124;
      end
      11'b00001111101 : begin
        result = input_125;
      end
      11'b00001111110 : begin
        result = input_126;
      end
      11'b00001111111 : begin
        result = input_127;
      end
      11'b00010000000 : begin
        result = input_128;
      end
      11'b00010000001 : begin
        result = input_129;
      end
      11'b00010000010 : begin
        result = input_130;
      end
      11'b00010000011 : begin
        result = input_131;
      end
      11'b00010000100 : begin
        result = input_132;
      end
      11'b00010000101 : begin
        result = input_133;
      end
      11'b00010000110 : begin
        result = input_134;
      end
      11'b00010000111 : begin
        result = input_135;
      end
      11'b00010001000 : begin
        result = input_136;
      end
      11'b00010001001 : begin
        result = input_137;
      end
      11'b00010001010 : begin
        result = input_138;
      end
      11'b00010001011 : begin
        result = input_139;
      end
      11'b00010001100 : begin
        result = input_140;
      end
      11'b00010001101 : begin
        result = input_141;
      end
      11'b00010001110 : begin
        result = input_142;
      end
      11'b00010001111 : begin
        result = input_143;
      end
      11'b00010010000 : begin
        result = input_144;
      end
      11'b00010010001 : begin
        result = input_145;
      end
      11'b00010010010 : begin
        result = input_146;
      end
      11'b00010010011 : begin
        result = input_147;
      end
      11'b00010010100 : begin
        result = input_148;
      end
      11'b00010010101 : begin
        result = input_149;
      end
      11'b00010010110 : begin
        result = input_150;
      end
      11'b00010010111 : begin
        result = input_151;
      end
      11'b00010011000 : begin
        result = input_152;
      end
      11'b00010011001 : begin
        result = input_153;
      end
      11'b00010011010 : begin
        result = input_154;
      end
      11'b00010011011 : begin
        result = input_155;
      end
      11'b00010011100 : begin
        result = input_156;
      end
      11'b00010011101 : begin
        result = input_157;
      end
      11'b00010011110 : begin
        result = input_158;
      end
      11'b00010011111 : begin
        result = input_159;
      end
      11'b00010100000 : begin
        result = input_160;
      end
      11'b00010100001 : begin
        result = input_161;
      end
      11'b00010100010 : begin
        result = input_162;
      end
      11'b00010100011 : begin
        result = input_163;
      end
      11'b00010100100 : begin
        result = input_164;
      end
      11'b00010100101 : begin
        result = input_165;
      end
      11'b00010100110 : begin
        result = input_166;
      end
      11'b00010100111 : begin
        result = input_167;
      end
      11'b00010101000 : begin
        result = input_168;
      end
      11'b00010101001 : begin
        result = input_169;
      end
      11'b00010101010 : begin
        result = input_170;
      end
      11'b00010101011 : begin
        result = input_171;
      end
      11'b00010101100 : begin
        result = input_172;
      end
      11'b00010101101 : begin
        result = input_173;
      end
      11'b00010101110 : begin
        result = input_174;
      end
      11'b00010101111 : begin
        result = input_175;
      end
      11'b00010110000 : begin
        result = input_176;
      end
      11'b00010110001 : begin
        result = input_177;
      end
      11'b00010110010 : begin
        result = input_178;
      end
      11'b00010110011 : begin
        result = input_179;
      end
      11'b00010110100 : begin
        result = input_180;
      end
      11'b00010110101 : begin
        result = input_181;
      end
      11'b00010110110 : begin
        result = input_182;
      end
      11'b00010110111 : begin
        result = input_183;
      end
      11'b00010111000 : begin
        result = input_184;
      end
      11'b00010111001 : begin
        result = input_185;
      end
      11'b00010111010 : begin
        result = input_186;
      end
      11'b00010111011 : begin
        result = input_187;
      end
      11'b00010111100 : begin
        result = input_188;
      end
      11'b00010111101 : begin
        result = input_189;
      end
      11'b00010111110 : begin
        result = input_190;
      end
      11'b00010111111 : begin
        result = input_191;
      end
      11'b00011000000 : begin
        result = input_192;
      end
      11'b00011000001 : begin
        result = input_193;
      end
      11'b00011000010 : begin
        result = input_194;
      end
      11'b00011000011 : begin
        result = input_195;
      end
      11'b00011000100 : begin
        result = input_196;
      end
      11'b00011000101 : begin
        result = input_197;
      end
      11'b00011000110 : begin
        result = input_198;
      end
      11'b00011000111 : begin
        result = input_199;
      end
      11'b00011001000 : begin
        result = input_200;
      end
      11'b00011001001 : begin
        result = input_201;
      end
      11'b00011001010 : begin
        result = input_202;
      end
      11'b00011001011 : begin
        result = input_203;
      end
      11'b00011001100 : begin
        result = input_204;
      end
      11'b00011001101 : begin
        result = input_205;
      end
      11'b00011001110 : begin
        result = input_206;
      end
      11'b00011001111 : begin
        result = input_207;
      end
      11'b00011010000 : begin
        result = input_208;
      end
      11'b00011010001 : begin
        result = input_209;
      end
      11'b00011010010 : begin
        result = input_210;
      end
      11'b00011010011 : begin
        result = input_211;
      end
      11'b00011010100 : begin
        result = input_212;
      end
      11'b00011010101 : begin
        result = input_213;
      end
      11'b00011010110 : begin
        result = input_214;
      end
      11'b00011010111 : begin
        result = input_215;
      end
      11'b00011011000 : begin
        result = input_216;
      end
      11'b00011011001 : begin
        result = input_217;
      end
      11'b00011011010 : begin
        result = input_218;
      end
      11'b00011011011 : begin
        result = input_219;
      end
      11'b00011011100 : begin
        result = input_220;
      end
      11'b00011011101 : begin
        result = input_221;
      end
      11'b00011011110 : begin
        result = input_222;
      end
      11'b00011011111 : begin
        result = input_223;
      end
      11'b00011100000 : begin
        result = input_224;
      end
      11'b00011100001 : begin
        result = input_225;
      end
      11'b00011100010 : begin
        result = input_226;
      end
      11'b00011100011 : begin
        result = input_227;
      end
      11'b00011100100 : begin
        result = input_228;
      end
      11'b00011100101 : begin
        result = input_229;
      end
      11'b00011100110 : begin
        result = input_230;
      end
      11'b00011100111 : begin
        result = input_231;
      end
      11'b00011101000 : begin
        result = input_232;
      end
      11'b00011101001 : begin
        result = input_233;
      end
      11'b00011101010 : begin
        result = input_234;
      end
      11'b00011101011 : begin
        result = input_235;
      end
      11'b00011101100 : begin
        result = input_236;
      end
      11'b00011101101 : begin
        result = input_237;
      end
      11'b00011101110 : begin
        result = input_238;
      end
      11'b00011101111 : begin
        result = input_239;
      end
      11'b00011110000 : begin
        result = input_240;
      end
      11'b00011110001 : begin
        result = input_241;
      end
      11'b00011110010 : begin
        result = input_242;
      end
      11'b00011110011 : begin
        result = input_243;
      end
      11'b00011110100 : begin
        result = input_244;
      end
      11'b00011110101 : begin
        result = input_245;
      end
      11'b00011110110 : begin
        result = input_246;
      end
      11'b00011110111 : begin
        result = input_247;
      end
      11'b00011111000 : begin
        result = input_248;
      end
      11'b00011111001 : begin
        result = input_249;
      end
      11'b00011111010 : begin
        result = input_250;
      end
      11'b00011111011 : begin
        result = input_251;
      end
      11'b00011111100 : begin
        result = input_252;
      end
      11'b00011111101 : begin
        result = input_253;
      end
      11'b00011111110 : begin
        result = input_254;
      end
      11'b00011111111 : begin
        result = input_255;
      end
      11'b00100000000 : begin
        result = input_256;
      end
      11'b00100000001 : begin
        result = input_257;
      end
      11'b00100000010 : begin
        result = input_258;
      end
      11'b00100000011 : begin
        result = input_259;
      end
      11'b00100000100 : begin
        result = input_260;
      end
      11'b00100000101 : begin
        result = input_261;
      end
      11'b00100000110 : begin
        result = input_262;
      end
      11'b00100000111 : begin
        result = input_263;
      end
      11'b00100001000 : begin
        result = input_264;
      end
      11'b00100001001 : begin
        result = input_265;
      end
      11'b00100001010 : begin
        result = input_266;
      end
      11'b00100001011 : begin
        result = input_267;
      end
      11'b00100001100 : begin
        result = input_268;
      end
      11'b00100001101 : begin
        result = input_269;
      end
      11'b00100001110 : begin
        result = input_270;
      end
      11'b00100001111 : begin
        result = input_271;
      end
      11'b00100010000 : begin
        result = input_272;
      end
      11'b00100010001 : begin
        result = input_273;
      end
      11'b00100010010 : begin
        result = input_274;
      end
      11'b00100010011 : begin
        result = input_275;
      end
      11'b00100010100 : begin
        result = input_276;
      end
      11'b00100010101 : begin
        result = input_277;
      end
      11'b00100010110 : begin
        result = input_278;
      end
      11'b00100010111 : begin
        result = input_279;
      end
      11'b00100011000 : begin
        result = input_280;
      end
      11'b00100011001 : begin
        result = input_281;
      end
      11'b00100011010 : begin
        result = input_282;
      end
      11'b00100011011 : begin
        result = input_283;
      end
      11'b00100011100 : begin
        result = input_284;
      end
      11'b00100011101 : begin
        result = input_285;
      end
      11'b00100011110 : begin
        result = input_286;
      end
      11'b00100011111 : begin
        result = input_287;
      end
      11'b00100100000 : begin
        result = input_288;
      end
      11'b00100100001 : begin
        result = input_289;
      end
      11'b00100100010 : begin
        result = input_290;
      end
      11'b00100100011 : begin
        result = input_291;
      end
      11'b00100100100 : begin
        result = input_292;
      end
      11'b00100100101 : begin
        result = input_293;
      end
      11'b00100100110 : begin
        result = input_294;
      end
      11'b00100100111 : begin
        result = input_295;
      end
      11'b00100101000 : begin
        result = input_296;
      end
      11'b00100101001 : begin
        result = input_297;
      end
      11'b00100101010 : begin
        result = input_298;
      end
      11'b00100101011 : begin
        result = input_299;
      end
      11'b00100101100 : begin
        result = input_300;
      end
      11'b00100101101 : begin
        result = input_301;
      end
      11'b00100101110 : begin
        result = input_302;
      end
      11'b00100101111 : begin
        result = input_303;
      end
      11'b00100110000 : begin
        result = input_304;
      end
      11'b00100110001 : begin
        result = input_305;
      end
      11'b00100110010 : begin
        result = input_306;
      end
      11'b00100110011 : begin
        result = input_307;
      end
      11'b00100110100 : begin
        result = input_308;
      end
      11'b00100110101 : begin
        result = input_309;
      end
      11'b00100110110 : begin
        result = input_310;
      end
      11'b00100110111 : begin
        result = input_311;
      end
      11'b00100111000 : begin
        result = input_312;
      end
      11'b00100111001 : begin
        result = input_313;
      end
      11'b00100111010 : begin
        result = input_314;
      end
      11'b00100111011 : begin
        result = input_315;
      end
      11'b00100111100 : begin
        result = input_316;
      end
      11'b00100111101 : begin
        result = input_317;
      end
      11'b00100111110 : begin
        result = input_318;
      end
      11'b00100111111 : begin
        result = input_319;
      end
      11'b00101000000 : begin
        result = input_320;
      end
      11'b00101000001 : begin
        result = input_321;
      end
      11'b00101000010 : begin
        result = input_322;
      end
      11'b00101000011 : begin
        result = input_323;
      end
      11'b00101000100 : begin
        result = input_324;
      end
      11'b00101000101 : begin
        result = input_325;
      end
      11'b00101000110 : begin
        result = input_326;
      end
      11'b00101000111 : begin
        result = input_327;
      end
      11'b00101001000 : begin
        result = input_328;
      end
      11'b00101001001 : begin
        result = input_329;
      end
      11'b00101001010 : begin
        result = input_330;
      end
      11'b00101001011 : begin
        result = input_331;
      end
      11'b00101001100 : begin
        result = input_332;
      end
      11'b00101001101 : begin
        result = input_333;
      end
      11'b00101001110 : begin
        result = input_334;
      end
      11'b00101001111 : begin
        result = input_335;
      end
      11'b00101010000 : begin
        result = input_336;
      end
      11'b00101010001 : begin
        result = input_337;
      end
      11'b00101010010 : begin
        result = input_338;
      end
      11'b00101010011 : begin
        result = input_339;
      end
      11'b00101010100 : begin
        result = input_340;
      end
      11'b00101010101 : begin
        result = input_341;
      end
      11'b00101010110 : begin
        result = input_342;
      end
      11'b00101010111 : begin
        result = input_343;
      end
      11'b00101011000 : begin
        result = input_344;
      end
      11'b00101011001 : begin
        result = input_345;
      end
      11'b00101011010 : begin
        result = input_346;
      end
      11'b00101011011 : begin
        result = input_347;
      end
      11'b00101011100 : begin
        result = input_348;
      end
      11'b00101011101 : begin
        result = input_349;
      end
      11'b00101011110 : begin
        result = input_350;
      end
      11'b00101011111 : begin
        result = input_351;
      end
      11'b00101100000 : begin
        result = input_352;
      end
      11'b00101100001 : begin
        result = input_353;
      end
      11'b00101100010 : begin
        result = input_354;
      end
      11'b00101100011 : begin
        result = input_355;
      end
      11'b00101100100 : begin
        result = input_356;
      end
      11'b00101100101 : begin
        result = input_357;
      end
      11'b00101100110 : begin
        result = input_358;
      end
      11'b00101100111 : begin
        result = input_359;
      end
      11'b00101101000 : begin
        result = input_360;
      end
      11'b00101101001 : begin
        result = input_361;
      end
      11'b00101101010 : begin
        result = input_362;
      end
      11'b00101101011 : begin
        result = input_363;
      end
      11'b00101101100 : begin
        result = input_364;
      end
      11'b00101101101 : begin
        result = input_365;
      end
      11'b00101101110 : begin
        result = input_366;
      end
      11'b00101101111 : begin
        result = input_367;
      end
      11'b00101110000 : begin
        result = input_368;
      end
      11'b00101110001 : begin
        result = input_369;
      end
      11'b00101110010 : begin
        result = input_370;
      end
      11'b00101110011 : begin
        result = input_371;
      end
      11'b00101110100 : begin
        result = input_372;
      end
      11'b00101110101 : begin
        result = input_373;
      end
      11'b00101110110 : begin
        result = input_374;
      end
      11'b00101110111 : begin
        result = input_375;
      end
      11'b00101111000 : begin
        result = input_376;
      end
      11'b00101111001 : begin
        result = input_377;
      end
      11'b00101111010 : begin
        result = input_378;
      end
      11'b00101111011 : begin
        result = input_379;
      end
      11'b00101111100 : begin
        result = input_380;
      end
      11'b00101111101 : begin
        result = input_381;
      end
      11'b00101111110 : begin
        result = input_382;
      end
      11'b00101111111 : begin
        result = input_383;
      end
      11'b00110000000 : begin
        result = input_384;
      end
      11'b00110000001 : begin
        result = input_385;
      end
      11'b00110000010 : begin
        result = input_386;
      end
      11'b00110000011 : begin
        result = input_387;
      end
      11'b00110000100 : begin
        result = input_388;
      end
      11'b00110000101 : begin
        result = input_389;
      end
      11'b00110000110 : begin
        result = input_390;
      end
      11'b00110000111 : begin
        result = input_391;
      end
      11'b00110001000 : begin
        result = input_392;
      end
      11'b00110001001 : begin
        result = input_393;
      end
      11'b00110001010 : begin
        result = input_394;
      end
      11'b00110001011 : begin
        result = input_395;
      end
      11'b00110001100 : begin
        result = input_396;
      end
      11'b00110001101 : begin
        result = input_397;
      end
      11'b00110001110 : begin
        result = input_398;
      end
      11'b00110001111 : begin
        result = input_399;
      end
      11'b00110010000 : begin
        result = input_400;
      end
      11'b00110010001 : begin
        result = input_401;
      end
      11'b00110010010 : begin
        result = input_402;
      end
      11'b00110010011 : begin
        result = input_403;
      end
      11'b00110010100 : begin
        result = input_404;
      end
      11'b00110010101 : begin
        result = input_405;
      end
      11'b00110010110 : begin
        result = input_406;
      end
      11'b00110010111 : begin
        result = input_407;
      end
      11'b00110011000 : begin
        result = input_408;
      end
      11'b00110011001 : begin
        result = input_409;
      end
      11'b00110011010 : begin
        result = input_410;
      end
      11'b00110011011 : begin
        result = input_411;
      end
      11'b00110011100 : begin
        result = input_412;
      end
      11'b00110011101 : begin
        result = input_413;
      end
      11'b00110011110 : begin
        result = input_414;
      end
      11'b00110011111 : begin
        result = input_415;
      end
      11'b00110100000 : begin
        result = input_416;
      end
      11'b00110100001 : begin
        result = input_417;
      end
      11'b00110100010 : begin
        result = input_418;
      end
      11'b00110100011 : begin
        result = input_419;
      end
      11'b00110100100 : begin
        result = input_420;
      end
      11'b00110100101 : begin
        result = input_421;
      end
      11'b00110100110 : begin
        result = input_422;
      end
      11'b00110100111 : begin
        result = input_423;
      end
      11'b00110101000 : begin
        result = input_424;
      end
      11'b00110101001 : begin
        result = input_425;
      end
      11'b00110101010 : begin
        result = input_426;
      end
      11'b00110101011 : begin
        result = input_427;
      end
      11'b00110101100 : begin
        result = input_428;
      end
      11'b00110101101 : begin
        result = input_429;
      end
      11'b00110101110 : begin
        result = input_430;
      end
      11'b00110101111 : begin
        result = input_431;
      end
      11'b00110110000 : begin
        result = input_432;
      end
      11'b00110110001 : begin
        result = input_433;
      end
      11'b00110110010 : begin
        result = input_434;
      end
      11'b00110110011 : begin
        result = input_435;
      end
      11'b00110110100 : begin
        result = input_436;
      end
      11'b00110110101 : begin
        result = input_437;
      end
      11'b00110110110 : begin
        result = input_438;
      end
      11'b00110110111 : begin
        result = input_439;
      end
      11'b00110111000 : begin
        result = input_440;
      end
      11'b00110111001 : begin
        result = input_441;
      end
      11'b00110111010 : begin
        result = input_442;
      end
      11'b00110111011 : begin
        result = input_443;
      end
      11'b00110111100 : begin
        result = input_444;
      end
      11'b00110111101 : begin
        result = input_445;
      end
      11'b00110111110 : begin
        result = input_446;
      end
      11'b00110111111 : begin
        result = input_447;
      end
      11'b00111000000 : begin
        result = input_448;
      end
      11'b00111000001 : begin
        result = input_449;
      end
      11'b00111000010 : begin
        result = input_450;
      end
      11'b00111000011 : begin
        result = input_451;
      end
      11'b00111000100 : begin
        result = input_452;
      end
      11'b00111000101 : begin
        result = input_453;
      end
      11'b00111000110 : begin
        result = input_454;
      end
      11'b00111000111 : begin
        result = input_455;
      end
      11'b00111001000 : begin
        result = input_456;
      end
      11'b00111001001 : begin
        result = input_457;
      end
      11'b00111001010 : begin
        result = input_458;
      end
      11'b00111001011 : begin
        result = input_459;
      end
      11'b00111001100 : begin
        result = input_460;
      end
      11'b00111001101 : begin
        result = input_461;
      end
      11'b00111001110 : begin
        result = input_462;
      end
      11'b00111001111 : begin
        result = input_463;
      end
      11'b00111010000 : begin
        result = input_464;
      end
      11'b00111010001 : begin
        result = input_465;
      end
      11'b00111010010 : begin
        result = input_466;
      end
      11'b00111010011 : begin
        result = input_467;
      end
      11'b00111010100 : begin
        result = input_468;
      end
      11'b00111010101 : begin
        result = input_469;
      end
      11'b00111010110 : begin
        result = input_470;
      end
      11'b00111010111 : begin
        result = input_471;
      end
      11'b00111011000 : begin
        result = input_472;
      end
      11'b00111011001 : begin
        result = input_473;
      end
      11'b00111011010 : begin
        result = input_474;
      end
      11'b00111011011 : begin
        result = input_475;
      end
      11'b00111011100 : begin
        result = input_476;
      end
      11'b00111011101 : begin
        result = input_477;
      end
      11'b00111011110 : begin
        result = input_478;
      end
      11'b00111011111 : begin
        result = input_479;
      end
      11'b00111100000 : begin
        result = input_480;
      end
      11'b00111100001 : begin
        result = input_481;
      end
      11'b00111100010 : begin
        result = input_482;
      end
      11'b00111100011 : begin
        result = input_483;
      end
      11'b00111100100 : begin
        result = input_484;
      end
      11'b00111100101 : begin
        result = input_485;
      end
      11'b00111100110 : begin
        result = input_486;
      end
      11'b00111100111 : begin
        result = input_487;
      end
      11'b00111101000 : begin
        result = input_488;
      end
      11'b00111101001 : begin
        result = input_489;
      end
      11'b00111101010 : begin
        result = input_490;
      end
      11'b00111101011 : begin
        result = input_491;
      end
      11'b00111101100 : begin
        result = input_492;
      end
      11'b00111101101 : begin
        result = input_493;
      end
      11'b00111101110 : begin
        result = input_494;
      end
      11'b00111101111 : begin
        result = input_495;
      end
      11'b00111110000 : begin
        result = input_496;
      end
      11'b00111110001 : begin
        result = input_497;
      end
      11'b00111110010 : begin
        result = input_498;
      end
      11'b00111110011 : begin
        result = input_499;
      end
      11'b00111110100 : begin
        result = input_500;
      end
      11'b00111110101 : begin
        result = input_501;
      end
      11'b00111110110 : begin
        result = input_502;
      end
      11'b00111110111 : begin
        result = input_503;
      end
      11'b00111111000 : begin
        result = input_504;
      end
      11'b00111111001 : begin
        result = input_505;
      end
      11'b00111111010 : begin
        result = input_506;
      end
      11'b00111111011 : begin
        result = input_507;
      end
      11'b00111111100 : begin
        result = input_508;
      end
      11'b00111111101 : begin
        result = input_509;
      end
      11'b00111111110 : begin
        result = input_510;
      end
      11'b00111111111 : begin
        result = input_511;
      end
      11'b01000000000 : begin
        result = input_512;
      end
      11'b01000000001 : begin
        result = input_513;
      end
      11'b01000000010 : begin
        result = input_514;
      end
      11'b01000000011 : begin
        result = input_515;
      end
      11'b01000000100 : begin
        result = input_516;
      end
      11'b01000000101 : begin
        result = input_517;
      end
      11'b01000000110 : begin
        result = input_518;
      end
      11'b01000000111 : begin
        result = input_519;
      end
      11'b01000001000 : begin
        result = input_520;
      end
      11'b01000001001 : begin
        result = input_521;
      end
      11'b01000001010 : begin
        result = input_522;
      end
      11'b01000001011 : begin
        result = input_523;
      end
      11'b01000001100 : begin
        result = input_524;
      end
      11'b01000001101 : begin
        result = input_525;
      end
      11'b01000001110 : begin
        result = input_526;
      end
      11'b01000001111 : begin
        result = input_527;
      end
      11'b01000010000 : begin
        result = input_528;
      end
      11'b01000010001 : begin
        result = input_529;
      end
      11'b01000010010 : begin
        result = input_530;
      end
      11'b01000010011 : begin
        result = input_531;
      end
      11'b01000010100 : begin
        result = input_532;
      end
      11'b01000010101 : begin
        result = input_533;
      end
      11'b01000010110 : begin
        result = input_534;
      end
      11'b01000010111 : begin
        result = input_535;
      end
      11'b01000011000 : begin
        result = input_536;
      end
      11'b01000011001 : begin
        result = input_537;
      end
      11'b01000011010 : begin
        result = input_538;
      end
      11'b01000011011 : begin
        result = input_539;
      end
      11'b01000011100 : begin
        result = input_540;
      end
      11'b01000011101 : begin
        result = input_541;
      end
      11'b01000011110 : begin
        result = input_542;
      end
      11'b01000011111 : begin
        result = input_543;
      end
      11'b01000100000 : begin
        result = input_544;
      end
      11'b01000100001 : begin
        result = input_545;
      end
      11'b01000100010 : begin
        result = input_546;
      end
      11'b01000100011 : begin
        result = input_547;
      end
      11'b01000100100 : begin
        result = input_548;
      end
      11'b01000100101 : begin
        result = input_549;
      end
      11'b01000100110 : begin
        result = input_550;
      end
      11'b01000100111 : begin
        result = input_551;
      end
      11'b01000101000 : begin
        result = input_552;
      end
      11'b01000101001 : begin
        result = input_553;
      end
      11'b01000101010 : begin
        result = input_554;
      end
      11'b01000101011 : begin
        result = input_555;
      end
      11'b01000101100 : begin
        result = input_556;
      end
      11'b01000101101 : begin
        result = input_557;
      end
      11'b01000101110 : begin
        result = input_558;
      end
      11'b01000101111 : begin
        result = input_559;
      end
      11'b01000110000 : begin
        result = input_560;
      end
      11'b01000110001 : begin
        result = input_561;
      end
      11'b01000110010 : begin
        result = input_562;
      end
      11'b01000110011 : begin
        result = input_563;
      end
      11'b01000110100 : begin
        result = input_564;
      end
      11'b01000110101 : begin
        result = input_565;
      end
      11'b01000110110 : begin
        result = input_566;
      end
      11'b01000110111 : begin
        result = input_567;
      end
      11'b01000111000 : begin
        result = input_568;
      end
      11'b01000111001 : begin
        result = input_569;
      end
      11'b01000111010 : begin
        result = input_570;
      end
      11'b01000111011 : begin
        result = input_571;
      end
      11'b01000111100 : begin
        result = input_572;
      end
      11'b01000111101 : begin
        result = input_573;
      end
      11'b01000111110 : begin
        result = input_574;
      end
      11'b01000111111 : begin
        result = input_575;
      end
      11'b01001000000 : begin
        result = input_576;
      end
      11'b01001000001 : begin
        result = input_577;
      end
      11'b01001000010 : begin
        result = input_578;
      end
      11'b01001000011 : begin
        result = input_579;
      end
      11'b01001000100 : begin
        result = input_580;
      end
      11'b01001000101 : begin
        result = input_581;
      end
      11'b01001000110 : begin
        result = input_582;
      end
      11'b01001000111 : begin
        result = input_583;
      end
      11'b01001001000 : begin
        result = input_584;
      end
      11'b01001001001 : begin
        result = input_585;
      end
      11'b01001001010 : begin
        result = input_586;
      end
      11'b01001001011 : begin
        result = input_587;
      end
      11'b01001001100 : begin
        result = input_588;
      end
      11'b01001001101 : begin
        result = input_589;
      end
      11'b01001001110 : begin
        result = input_590;
      end
      11'b01001001111 : begin
        result = input_591;
      end
      11'b01001010000 : begin
        result = input_592;
      end
      11'b01001010001 : begin
        result = input_593;
      end
      11'b01001010010 : begin
        result = input_594;
      end
      11'b01001010011 : begin
        result = input_595;
      end
      11'b01001010100 : begin
        result = input_596;
      end
      11'b01001010101 : begin
        result = input_597;
      end
      11'b01001010110 : begin
        result = input_598;
      end
      11'b01001010111 : begin
        result = input_599;
      end
      11'b01001011000 : begin
        result = input_600;
      end
      11'b01001011001 : begin
        result = input_601;
      end
      11'b01001011010 : begin
        result = input_602;
      end
      11'b01001011011 : begin
        result = input_603;
      end
      11'b01001011100 : begin
        result = input_604;
      end
      11'b01001011101 : begin
        result = input_605;
      end
      11'b01001011110 : begin
        result = input_606;
      end
      11'b01001011111 : begin
        result = input_607;
      end
      11'b01001100000 : begin
        result = input_608;
      end
      11'b01001100001 : begin
        result = input_609;
      end
      11'b01001100010 : begin
        result = input_610;
      end
      11'b01001100011 : begin
        result = input_611;
      end
      11'b01001100100 : begin
        result = input_612;
      end
      11'b01001100101 : begin
        result = input_613;
      end
      11'b01001100110 : begin
        result = input_614;
      end
      11'b01001100111 : begin
        result = input_615;
      end
      11'b01001101000 : begin
        result = input_616;
      end
      11'b01001101001 : begin
        result = input_617;
      end
      11'b01001101010 : begin
        result = input_618;
      end
      11'b01001101011 : begin
        result = input_619;
      end
      11'b01001101100 : begin
        result = input_620;
      end
      11'b01001101101 : begin
        result = input_621;
      end
      11'b01001101110 : begin
        result = input_622;
      end
      11'b01001101111 : begin
        result = input_623;
      end
      11'b01001110000 : begin
        result = input_624;
      end
      11'b01001110001 : begin
        result = input_625;
      end
      11'b01001110010 : begin
        result = input_626;
      end
      11'b01001110011 : begin
        result = input_627;
      end
      11'b01001110100 : begin
        result = input_628;
      end
      11'b01001110101 : begin
        result = input_629;
      end
      11'b01001110110 : begin
        result = input_630;
      end
      11'b01001110111 : begin
        result = input_631;
      end
      11'b01001111000 : begin
        result = input_632;
      end
      11'b01001111001 : begin
        result = input_633;
      end
      11'b01001111010 : begin
        result = input_634;
      end
      11'b01001111011 : begin
        result = input_635;
      end
      11'b01001111100 : begin
        result = input_636;
      end
      11'b01001111101 : begin
        result = input_637;
      end
      11'b01001111110 : begin
        result = input_638;
      end
      11'b01001111111 : begin
        result = input_639;
      end
      11'b01010000000 : begin
        result = input_640;
      end
      11'b01010000001 : begin
        result = input_641;
      end
      11'b01010000010 : begin
        result = input_642;
      end
      11'b01010000011 : begin
        result = input_643;
      end
      11'b01010000100 : begin
        result = input_644;
      end
      11'b01010000101 : begin
        result = input_645;
      end
      11'b01010000110 : begin
        result = input_646;
      end
      11'b01010000111 : begin
        result = input_647;
      end
      11'b01010001000 : begin
        result = input_648;
      end
      11'b01010001001 : begin
        result = input_649;
      end
      11'b01010001010 : begin
        result = input_650;
      end
      11'b01010001011 : begin
        result = input_651;
      end
      11'b01010001100 : begin
        result = input_652;
      end
      11'b01010001101 : begin
        result = input_653;
      end
      11'b01010001110 : begin
        result = input_654;
      end
      11'b01010001111 : begin
        result = input_655;
      end
      11'b01010010000 : begin
        result = input_656;
      end
      11'b01010010001 : begin
        result = input_657;
      end
      11'b01010010010 : begin
        result = input_658;
      end
      11'b01010010011 : begin
        result = input_659;
      end
      11'b01010010100 : begin
        result = input_660;
      end
      11'b01010010101 : begin
        result = input_661;
      end
      11'b01010010110 : begin
        result = input_662;
      end
      11'b01010010111 : begin
        result = input_663;
      end
      11'b01010011000 : begin
        result = input_664;
      end
      11'b01010011001 : begin
        result = input_665;
      end
      11'b01010011010 : begin
        result = input_666;
      end
      11'b01010011011 : begin
        result = input_667;
      end
      11'b01010011100 : begin
        result = input_668;
      end
      11'b01010011101 : begin
        result = input_669;
      end
      11'b01010011110 : begin
        result = input_670;
      end
      11'b01010011111 : begin
        result = input_671;
      end
      11'b01010100000 : begin
        result = input_672;
      end
      11'b01010100001 : begin
        result = input_673;
      end
      11'b01010100010 : begin
        result = input_674;
      end
      11'b01010100011 : begin
        result = input_675;
      end
      11'b01010100100 : begin
        result = input_676;
      end
      11'b01010100101 : begin
        result = input_677;
      end
      11'b01010100110 : begin
        result = input_678;
      end
      11'b01010100111 : begin
        result = input_679;
      end
      11'b01010101000 : begin
        result = input_680;
      end
      11'b01010101001 : begin
        result = input_681;
      end
      11'b01010101010 : begin
        result = input_682;
      end
      11'b01010101011 : begin
        result = input_683;
      end
      11'b01010101100 : begin
        result = input_684;
      end
      11'b01010101101 : begin
        result = input_685;
      end
      11'b01010101110 : begin
        result = input_686;
      end
      11'b01010101111 : begin
        result = input_687;
      end
      11'b01010110000 : begin
        result = input_688;
      end
      11'b01010110001 : begin
        result = input_689;
      end
      11'b01010110010 : begin
        result = input_690;
      end
      11'b01010110011 : begin
        result = input_691;
      end
      11'b01010110100 : begin
        result = input_692;
      end
      11'b01010110101 : begin
        result = input_693;
      end
      11'b01010110110 : begin
        result = input_694;
      end
      11'b01010110111 : begin
        result = input_695;
      end
      11'b01010111000 : begin
        result = input_696;
      end
      11'b01010111001 : begin
        result = input_697;
      end
      11'b01010111010 : begin
        result = input_698;
      end
      11'b01010111011 : begin
        result = input_699;
      end
      11'b01010111100 : begin
        result = input_700;
      end
      11'b01010111101 : begin
        result = input_701;
      end
      11'b01010111110 : begin
        result = input_702;
      end
      11'b01010111111 : begin
        result = input_703;
      end
      11'b01011000000 : begin
        result = input_704;
      end
      11'b01011000001 : begin
        result = input_705;
      end
      11'b01011000010 : begin
        result = input_706;
      end
      11'b01011000011 : begin
        result = input_707;
      end
      11'b01011000100 : begin
        result = input_708;
      end
      11'b01011000101 : begin
        result = input_709;
      end
      11'b01011000110 : begin
        result = input_710;
      end
      11'b01011000111 : begin
        result = input_711;
      end
      11'b01011001000 : begin
        result = input_712;
      end
      11'b01011001001 : begin
        result = input_713;
      end
      11'b01011001010 : begin
        result = input_714;
      end
      11'b01011001011 : begin
        result = input_715;
      end
      11'b01011001100 : begin
        result = input_716;
      end
      11'b01011001101 : begin
        result = input_717;
      end
      11'b01011001110 : begin
        result = input_718;
      end
      11'b01011001111 : begin
        result = input_719;
      end
      11'b01011010000 : begin
        result = input_720;
      end
      11'b01011010001 : begin
        result = input_721;
      end
      11'b01011010010 : begin
        result = input_722;
      end
      11'b01011010011 : begin
        result = input_723;
      end
      11'b01011010100 : begin
        result = input_724;
      end
      11'b01011010101 : begin
        result = input_725;
      end
      11'b01011010110 : begin
        result = input_726;
      end
      11'b01011010111 : begin
        result = input_727;
      end
      11'b01011011000 : begin
        result = input_728;
      end
      11'b01011011001 : begin
        result = input_729;
      end
      11'b01011011010 : begin
        result = input_730;
      end
      11'b01011011011 : begin
        result = input_731;
      end
      11'b01011011100 : begin
        result = input_732;
      end
      11'b01011011101 : begin
        result = input_733;
      end
      11'b01011011110 : begin
        result = input_734;
      end
      11'b01011011111 : begin
        result = input_735;
      end
      11'b01011100000 : begin
        result = input_736;
      end
      11'b01011100001 : begin
        result = input_737;
      end
      11'b01011100010 : begin
        result = input_738;
      end
      11'b01011100011 : begin
        result = input_739;
      end
      11'b01011100100 : begin
        result = input_740;
      end
      11'b01011100101 : begin
        result = input_741;
      end
      11'b01011100110 : begin
        result = input_742;
      end
      11'b01011100111 : begin
        result = input_743;
      end
      11'b01011101000 : begin
        result = input_744;
      end
      11'b01011101001 : begin
        result = input_745;
      end
      11'b01011101010 : begin
        result = input_746;
      end
      11'b01011101011 : begin
        result = input_747;
      end
      11'b01011101100 : begin
        result = input_748;
      end
      11'b01011101101 : begin
        result = input_749;
      end
      11'b01011101110 : begin
        result = input_750;
      end
      11'b01011101111 : begin
        result = input_751;
      end
      11'b01011110000 : begin
        result = input_752;
      end
      11'b01011110001 : begin
        result = input_753;
      end
      11'b01011110010 : begin
        result = input_754;
      end
      11'b01011110011 : begin
        result = input_755;
      end
      11'b01011110100 : begin
        result = input_756;
      end
      11'b01011110101 : begin
        result = input_757;
      end
      11'b01011110110 : begin
        result = input_758;
      end
      11'b01011110111 : begin
        result = input_759;
      end
      11'b01011111000 : begin
        result = input_760;
      end
      11'b01011111001 : begin
        result = input_761;
      end
      11'b01011111010 : begin
        result = input_762;
      end
      11'b01011111011 : begin
        result = input_763;
      end
      11'b01011111100 : begin
        result = input_764;
      end
      11'b01011111101 : begin
        result = input_765;
      end
      11'b01011111110 : begin
        result = input_766;
      end
      11'b01011111111 : begin
        result = input_767;
      end
      11'b01100000000 : begin
        result = input_768;
      end
      11'b01100000001 : begin
        result = input_769;
      end
      11'b01100000010 : begin
        result = input_770;
      end
      11'b01100000011 : begin
        result = input_771;
      end
      11'b01100000100 : begin
        result = input_772;
      end
      11'b01100000101 : begin
        result = input_773;
      end
      11'b01100000110 : begin
        result = input_774;
      end
      11'b01100000111 : begin
        result = input_775;
      end
      11'b01100001000 : begin
        result = input_776;
      end
      11'b01100001001 : begin
        result = input_777;
      end
      11'b01100001010 : begin
        result = input_778;
      end
      11'b01100001011 : begin
        result = input_779;
      end
      11'b01100001100 : begin
        result = input_780;
      end
      11'b01100001101 : begin
        result = input_781;
      end
      11'b01100001110 : begin
        result = input_782;
      end
      11'b01100001111 : begin
        result = input_783;
      end
      11'b01100010000 : begin
        result = input_784;
      end
      11'b01100010001 : begin
        result = input_785;
      end
      11'b01100010010 : begin
        result = input_786;
      end
      11'b01100010011 : begin
        result = input_787;
      end
      11'b01100010100 : begin
        result = input_788;
      end
      11'b01100010101 : begin
        result = input_789;
      end
      11'b01100010110 : begin
        result = input_790;
      end
      11'b01100010111 : begin
        result = input_791;
      end
      11'b01100011000 : begin
        result = input_792;
      end
      11'b01100011001 : begin
        result = input_793;
      end
      11'b01100011010 : begin
        result = input_794;
      end
      11'b01100011011 : begin
        result = input_795;
      end
      11'b01100011100 : begin
        result = input_796;
      end
      11'b01100011101 : begin
        result = input_797;
      end
      11'b01100011110 : begin
        result = input_798;
      end
      11'b01100011111 : begin
        result = input_799;
      end
      11'b01100100000 : begin
        result = input_800;
      end
      11'b01100100001 : begin
        result = input_801;
      end
      11'b01100100010 : begin
        result = input_802;
      end
      11'b01100100011 : begin
        result = input_803;
      end
      11'b01100100100 : begin
        result = input_804;
      end
      11'b01100100101 : begin
        result = input_805;
      end
      11'b01100100110 : begin
        result = input_806;
      end
      11'b01100100111 : begin
        result = input_807;
      end
      11'b01100101000 : begin
        result = input_808;
      end
      11'b01100101001 : begin
        result = input_809;
      end
      11'b01100101010 : begin
        result = input_810;
      end
      11'b01100101011 : begin
        result = input_811;
      end
      11'b01100101100 : begin
        result = input_812;
      end
      11'b01100101101 : begin
        result = input_813;
      end
      11'b01100101110 : begin
        result = input_814;
      end
      11'b01100101111 : begin
        result = input_815;
      end
      11'b01100110000 : begin
        result = input_816;
      end
      11'b01100110001 : begin
        result = input_817;
      end
      11'b01100110010 : begin
        result = input_818;
      end
      11'b01100110011 : begin
        result = input_819;
      end
      11'b01100110100 : begin
        result = input_820;
      end
      11'b01100110101 : begin
        result = input_821;
      end
      11'b01100110110 : begin
        result = input_822;
      end
      11'b01100110111 : begin
        result = input_823;
      end
      11'b01100111000 : begin
        result = input_824;
      end
      11'b01100111001 : begin
        result = input_825;
      end
      11'b01100111010 : begin
        result = input_826;
      end
      11'b01100111011 : begin
        result = input_827;
      end
      11'b01100111100 : begin
        result = input_828;
      end
      11'b01100111101 : begin
        result = input_829;
      end
      11'b01100111110 : begin
        result = input_830;
      end
      11'b01100111111 : begin
        result = input_831;
      end
      11'b01101000000 : begin
        result = input_832;
      end
      11'b01101000001 : begin
        result = input_833;
      end
      11'b01101000010 : begin
        result = input_834;
      end
      11'b01101000011 : begin
        result = input_835;
      end
      11'b01101000100 : begin
        result = input_836;
      end
      11'b01101000101 : begin
        result = input_837;
      end
      11'b01101000110 : begin
        result = input_838;
      end
      11'b01101000111 : begin
        result = input_839;
      end
      11'b01101001000 : begin
        result = input_840;
      end
      11'b01101001001 : begin
        result = input_841;
      end
      11'b01101001010 : begin
        result = input_842;
      end
      11'b01101001011 : begin
        result = input_843;
      end
      11'b01101001100 : begin
        result = input_844;
      end
      11'b01101001101 : begin
        result = input_845;
      end
      11'b01101001110 : begin
        result = input_846;
      end
      11'b01101001111 : begin
        result = input_847;
      end
      11'b01101010000 : begin
        result = input_848;
      end
      11'b01101010001 : begin
        result = input_849;
      end
      11'b01101010010 : begin
        result = input_850;
      end
      11'b01101010011 : begin
        result = input_851;
      end
      11'b01101010100 : begin
        result = input_852;
      end
      11'b01101010101 : begin
        result = input_853;
      end
      11'b01101010110 : begin
        result = input_854;
      end
      11'b01101010111 : begin
        result = input_855;
      end
      11'b01101011000 : begin
        result = input_856;
      end
      11'b01101011001 : begin
        result = input_857;
      end
      11'b01101011010 : begin
        result = input_858;
      end
      11'b01101011011 : begin
        result = input_859;
      end
      11'b01101011100 : begin
        result = input_860;
      end
      11'b01101011101 : begin
        result = input_861;
      end
      11'b01101011110 : begin
        result = input_862;
      end
      11'b01101011111 : begin
        result = input_863;
      end
      11'b01101100000 : begin
        result = input_864;
      end
      11'b01101100001 : begin
        result = input_865;
      end
      11'b01101100010 : begin
        result = input_866;
      end
      11'b01101100011 : begin
        result = input_867;
      end
      11'b01101100100 : begin
        result = input_868;
      end
      11'b01101100101 : begin
        result = input_869;
      end
      11'b01101100110 : begin
        result = input_870;
      end
      11'b01101100111 : begin
        result = input_871;
      end
      11'b01101101000 : begin
        result = input_872;
      end
      11'b01101101001 : begin
        result = input_873;
      end
      11'b01101101010 : begin
        result = input_874;
      end
      11'b01101101011 : begin
        result = input_875;
      end
      11'b01101101100 : begin
        result = input_876;
      end
      11'b01101101101 : begin
        result = input_877;
      end
      11'b01101101110 : begin
        result = input_878;
      end
      11'b01101101111 : begin
        result = input_879;
      end
      11'b01101110000 : begin
        result = input_880;
      end
      11'b01101110001 : begin
        result = input_881;
      end
      11'b01101110010 : begin
        result = input_882;
      end
      11'b01101110011 : begin
        result = input_883;
      end
      11'b01101110100 : begin
        result = input_884;
      end
      11'b01101110101 : begin
        result = input_885;
      end
      11'b01101110110 : begin
        result = input_886;
      end
      11'b01101110111 : begin
        result = input_887;
      end
      11'b01101111000 : begin
        result = input_888;
      end
      11'b01101111001 : begin
        result = input_889;
      end
      11'b01101111010 : begin
        result = input_890;
      end
      11'b01101111011 : begin
        result = input_891;
      end
      11'b01101111100 : begin
        result = input_892;
      end
      11'b01101111101 : begin
        result = input_893;
      end
      11'b01101111110 : begin
        result = input_894;
      end
      11'b01101111111 : begin
        result = input_895;
      end
      11'b01110000000 : begin
        result = input_896;
      end
      11'b01110000001 : begin
        result = input_897;
      end
      11'b01110000010 : begin
        result = input_898;
      end
      11'b01110000011 : begin
        result = input_899;
      end
      11'b01110000100 : begin
        result = input_900;
      end
      11'b01110000101 : begin
        result = input_901;
      end
      11'b01110000110 : begin
        result = input_902;
      end
      11'b01110000111 : begin
        result = input_903;
      end
      11'b01110001000 : begin
        result = input_904;
      end
      11'b01110001001 : begin
        result = input_905;
      end
      11'b01110001010 : begin
        result = input_906;
      end
      11'b01110001011 : begin
        result = input_907;
      end
      11'b01110001100 : begin
        result = input_908;
      end
      11'b01110001101 : begin
        result = input_909;
      end
      11'b01110001110 : begin
        result = input_910;
      end
      11'b01110001111 : begin
        result = input_911;
      end
      11'b01110010000 : begin
        result = input_912;
      end
      11'b01110010001 : begin
        result = input_913;
      end
      11'b01110010010 : begin
        result = input_914;
      end
      11'b01110010011 : begin
        result = input_915;
      end
      11'b01110010100 : begin
        result = input_916;
      end
      11'b01110010101 : begin
        result = input_917;
      end
      11'b01110010110 : begin
        result = input_918;
      end
      11'b01110010111 : begin
        result = input_919;
      end
      11'b01110011000 : begin
        result = input_920;
      end
      11'b01110011001 : begin
        result = input_921;
      end
      11'b01110011010 : begin
        result = input_922;
      end
      11'b01110011011 : begin
        result = input_923;
      end
      11'b01110011100 : begin
        result = input_924;
      end
      11'b01110011101 : begin
        result = input_925;
      end
      11'b01110011110 : begin
        result = input_926;
      end
      11'b01110011111 : begin
        result = input_927;
      end
      11'b01110100000 : begin
        result = input_928;
      end
      11'b01110100001 : begin
        result = input_929;
      end
      11'b01110100010 : begin
        result = input_930;
      end
      11'b01110100011 : begin
        result = input_931;
      end
      11'b01110100100 : begin
        result = input_932;
      end
      11'b01110100101 : begin
        result = input_933;
      end
      11'b01110100110 : begin
        result = input_934;
      end
      11'b01110100111 : begin
        result = input_935;
      end
      11'b01110101000 : begin
        result = input_936;
      end
      11'b01110101001 : begin
        result = input_937;
      end
      11'b01110101010 : begin
        result = input_938;
      end
      11'b01110101011 : begin
        result = input_939;
      end
      11'b01110101100 : begin
        result = input_940;
      end
      11'b01110101101 : begin
        result = input_941;
      end
      11'b01110101110 : begin
        result = input_942;
      end
      11'b01110101111 : begin
        result = input_943;
      end
      11'b01110110000 : begin
        result = input_944;
      end
      11'b01110110001 : begin
        result = input_945;
      end
      11'b01110110010 : begin
        result = input_946;
      end
      11'b01110110011 : begin
        result = input_947;
      end
      11'b01110110100 : begin
        result = input_948;
      end
      11'b01110110101 : begin
        result = input_949;
      end
      11'b01110110110 : begin
        result = input_950;
      end
      11'b01110110111 : begin
        result = input_951;
      end
      11'b01110111000 : begin
        result = input_952;
      end
      11'b01110111001 : begin
        result = input_953;
      end
      11'b01110111010 : begin
        result = input_954;
      end
      11'b01110111011 : begin
        result = input_955;
      end
      11'b01110111100 : begin
        result = input_956;
      end
      11'b01110111101 : begin
        result = input_957;
      end
      11'b01110111110 : begin
        result = input_958;
      end
      11'b01110111111 : begin
        result = input_959;
      end
      11'b01111000000 : begin
        result = input_960;
      end
      11'b01111000001 : begin
        result = input_961;
      end
      11'b01111000010 : begin
        result = input_962;
      end
      11'b01111000011 : begin
        result = input_963;
      end
      11'b01111000100 : begin
        result = input_964;
      end
      11'b01111000101 : begin
        result = input_965;
      end
      11'b01111000110 : begin
        result = input_966;
      end
      11'b01111000111 : begin
        result = input_967;
      end
      11'b01111001000 : begin
        result = input_968;
      end
      11'b01111001001 : begin
        result = input_969;
      end
      11'b01111001010 : begin
        result = input_970;
      end
      11'b01111001011 : begin
        result = input_971;
      end
      11'b01111001100 : begin
        result = input_972;
      end
      11'b01111001101 : begin
        result = input_973;
      end
      11'b01111001110 : begin
        result = input_974;
      end
      11'b01111001111 : begin
        result = input_975;
      end
      11'b01111010000 : begin
        result = input_976;
      end
      11'b01111010001 : begin
        result = input_977;
      end
      11'b01111010010 : begin
        result = input_978;
      end
      11'b01111010011 : begin
        result = input_979;
      end
      11'b01111010100 : begin
        result = input_980;
      end
      11'b01111010101 : begin
        result = input_981;
      end
      11'b01111010110 : begin
        result = input_982;
      end
      11'b01111010111 : begin
        result = input_983;
      end
      11'b01111011000 : begin
        result = input_984;
      end
      11'b01111011001 : begin
        result = input_985;
      end
      11'b01111011010 : begin
        result = input_986;
      end
      11'b01111011011 : begin
        result = input_987;
      end
      11'b01111011100 : begin
        result = input_988;
      end
      11'b01111011101 : begin
        result = input_989;
      end
      11'b01111011110 : begin
        result = input_990;
      end
      11'b01111011111 : begin
        result = input_991;
      end
      11'b01111100000 : begin
        result = input_992;
      end
      11'b01111100001 : begin
        result = input_993;
      end
      11'b01111100010 : begin
        result = input_994;
      end
      11'b01111100011 : begin
        result = input_995;
      end
      11'b01111100100 : begin
        result = input_996;
      end
      11'b01111100101 : begin
        result = input_997;
      end
      11'b01111100110 : begin
        result = input_998;
      end
      11'b01111100111 : begin
        result = input_999;
      end
      11'b01111101000 : begin
        result = input_1000;
      end
      11'b01111101001 : begin
        result = input_1001;
      end
      11'b01111101010 : begin
        result = input_1002;
      end
      11'b01111101011 : begin
        result = input_1003;
      end
      11'b01111101100 : begin
        result = input_1004;
      end
      11'b01111101101 : begin
        result = input_1005;
      end
      11'b01111101110 : begin
        result = input_1006;
      end
      11'b01111101111 : begin
        result = input_1007;
      end
      11'b01111110000 : begin
        result = input_1008;
      end
      11'b01111110001 : begin
        result = input_1009;
      end
      11'b01111110010 : begin
        result = input_1010;
      end
      11'b01111110011 : begin
        result = input_1011;
      end
      11'b01111110100 : begin
        result = input_1012;
      end
      11'b01111110101 : begin
        result = input_1013;
      end
      11'b01111110110 : begin
        result = input_1014;
      end
      11'b01111110111 : begin
        result = input_1015;
      end
      11'b01111111000 : begin
        result = input_1016;
      end
      11'b01111111001 : begin
        result = input_1017;
      end
      11'b01111111010 : begin
        result = input_1018;
      end
      11'b01111111011 : begin
        result = input_1019;
      end
      11'b01111111100 : begin
        result = input_1020;
      end
      11'b01111111101 : begin
        result = input_1021;
      end
      11'b01111111110 : begin
        result = input_1022;
      end
      11'b01111111111 : begin
        result = input_1023;
      end
      11'b10000000000 : begin
        result = input_1024;
      end
      11'b10000000001 : begin
        result = input_1025;
      end
      11'b10000000010 : begin
        result = input_1026;
      end
      11'b10000000011 : begin
        result = input_1027;
      end
      11'b10000000100 : begin
        result = input_1028;
      end
      11'b10000000101 : begin
        result = input_1029;
      end
      11'b10000000110 : begin
        result = input_1030;
      end
      11'b10000000111 : begin
        result = input_1031;
      end
      11'b10000001000 : begin
        result = input_1032;
      end
      11'b10000001001 : begin
        result = input_1033;
      end
      11'b10000001010 : begin
        result = input_1034;
      end
      11'b10000001011 : begin
        result = input_1035;
      end
      11'b10000001100 : begin
        result = input_1036;
      end
      11'b10000001101 : begin
        result = input_1037;
      end
      11'b10000001110 : begin
        result = input_1038;
      end
      11'b10000001111 : begin
        result = input_1039;
      end
      11'b10000010000 : begin
        result = input_1040;
      end
      11'b10000010001 : begin
        result = input_1041;
      end
      11'b10000010010 : begin
        result = input_1042;
      end
      11'b10000010011 : begin
        result = input_1043;
      end
      11'b10000010100 : begin
        result = input_1044;
      end
      11'b10000010101 : begin
        result = input_1045;
      end
      11'b10000010110 : begin
        result = input_1046;
      end
      11'b10000010111 : begin
        result = input_1047;
      end
      11'b10000011000 : begin
        result = input_1048;
      end
      11'b10000011001 : begin
        result = input_1049;
      end
      11'b10000011010 : begin
        result = input_1050;
      end
      11'b10000011011 : begin
        result = input_1051;
      end
      11'b10000011100 : begin
        result = input_1052;
      end
      11'b10000011101 : begin
        result = input_1053;
      end
      11'b10000011110 : begin
        result = input_1054;
      end
      11'b10000011111 : begin
        result = input_1055;
      end
      11'b10000100000 : begin
        result = input_1056;
      end
      11'b10000100001 : begin
        result = input_1057;
      end
      11'b10000100010 : begin
        result = input_1058;
      end
      11'b10000100011 : begin
        result = input_1059;
      end
      11'b10000100100 : begin
        result = input_1060;
      end
      11'b10000100101 : begin
        result = input_1061;
      end
      11'b10000100110 : begin
        result = input_1062;
      end
      11'b10000100111 : begin
        result = input_1063;
      end
      11'b10000101000 : begin
        result = input_1064;
      end
      11'b10000101001 : begin
        result = input_1065;
      end
      11'b10000101010 : begin
        result = input_1066;
      end
      11'b10000101011 : begin
        result = input_1067;
      end
      11'b10000101100 : begin
        result = input_1068;
      end
      11'b10000101101 : begin
        result = input_1069;
      end
      11'b10000101110 : begin
        result = input_1070;
      end
      11'b10000101111 : begin
        result = input_1071;
      end
      11'b10000110000 : begin
        result = input_1072;
      end
      11'b10000110001 : begin
        result = input_1073;
      end
      11'b10000110010 : begin
        result = input_1074;
      end
      11'b10000110011 : begin
        result = input_1075;
      end
      11'b10000110100 : begin
        result = input_1076;
      end
      11'b10000110101 : begin
        result = input_1077;
      end
      11'b10000110110 : begin
        result = input_1078;
      end
      11'b10000110111 : begin
        result = input_1079;
      end
      11'b10000111000 : begin
        result = input_1080;
      end
      11'b10000111001 : begin
        result = input_1081;
      end
      11'b10000111010 : begin
        result = input_1082;
      end
      11'b10000111011 : begin
        result = input_1083;
      end
      11'b10000111100 : begin
        result = input_1084;
      end
      11'b10000111101 : begin
        result = input_1085;
      end
      11'b10000111110 : begin
        result = input_1086;
      end
      11'b10000111111 : begin
        result = input_1087;
      end
      11'b10001000000 : begin
        result = input_1088;
      end
      11'b10001000001 : begin
        result = input_1089;
      end
      11'b10001000010 : begin
        result = input_1090;
      end
      11'b10001000011 : begin
        result = input_1091;
      end
      11'b10001000100 : begin
        result = input_1092;
      end
      11'b10001000101 : begin
        result = input_1093;
      end
      11'b10001000110 : begin
        result = input_1094;
      end
      11'b10001000111 : begin
        result = input_1095;
      end
      11'b10001001000 : begin
        result = input_1096;
      end
      11'b10001001001 : begin
        result = input_1097;
      end
      11'b10001001010 : begin
        result = input_1098;
      end
      11'b10001001011 : begin
        result = input_1099;
      end
      11'b10001001100 : begin
        result = input_1100;
      end
      11'b10001001101 : begin
        result = input_1101;
      end
      11'b10001001110 : begin
        result = input_1102;
      end
      11'b10001001111 : begin
        result = input_1103;
      end
      11'b10001010000 : begin
        result = input_1104;
      end
      11'b10001010001 : begin
        result = input_1105;
      end
      11'b10001010010 : begin
        result = input_1106;
      end
      11'b10001010011 : begin
        result = input_1107;
      end
      11'b10001010100 : begin
        result = input_1108;
      end
      11'b10001010101 : begin
        result = input_1109;
      end
      11'b10001010110 : begin
        result = input_1110;
      end
      11'b10001010111 : begin
        result = input_1111;
      end
      11'b10001011000 : begin
        result = input_1112;
      end
      11'b10001011001 : begin
        result = input_1113;
      end
      11'b10001011010 : begin
        result = input_1114;
      end
      11'b10001011011 : begin
        result = input_1115;
      end
      11'b10001011100 : begin
        result = input_1116;
      end
      11'b10001011101 : begin
        result = input_1117;
      end
      11'b10001011110 : begin
        result = input_1118;
      end
      11'b10001011111 : begin
        result = input_1119;
      end
      11'b10001100000 : begin
        result = input_1120;
      end
      11'b10001100001 : begin
        result = input_1121;
      end
      11'b10001100010 : begin
        result = input_1122;
      end
      11'b10001100011 : begin
        result = input_1123;
      end
      11'b10001100100 : begin
        result = input_1124;
      end
      11'b10001100101 : begin
        result = input_1125;
      end
      11'b10001100110 : begin
        result = input_1126;
      end
      11'b10001100111 : begin
        result = input_1127;
      end
      11'b10001101000 : begin
        result = input_1128;
      end
      11'b10001101001 : begin
        result = input_1129;
      end
      11'b10001101010 : begin
        result = input_1130;
      end
      11'b10001101011 : begin
        result = input_1131;
      end
      11'b10001101100 : begin
        result = input_1132;
      end
      11'b10001101101 : begin
        result = input_1133;
      end
      11'b10001101110 : begin
        result = input_1134;
      end
      11'b10001101111 : begin
        result = input_1135;
      end
      11'b10001110000 : begin
        result = input_1136;
      end
      11'b10001110001 : begin
        result = input_1137;
      end
      11'b10001110010 : begin
        result = input_1138;
      end
      11'b10001110011 : begin
        result = input_1139;
      end
      11'b10001110100 : begin
        result = input_1140;
      end
      11'b10001110101 : begin
        result = input_1141;
      end
      11'b10001110110 : begin
        result = input_1142;
      end
      11'b10001110111 : begin
        result = input_1143;
      end
      11'b10001111000 : begin
        result = input_1144;
      end
      11'b10001111001 : begin
        result = input_1145;
      end
      11'b10001111010 : begin
        result = input_1146;
      end
      11'b10001111011 : begin
        result = input_1147;
      end
      11'b10001111100 : begin
        result = input_1148;
      end
      11'b10001111101 : begin
        result = input_1149;
      end
      11'b10001111110 : begin
        result = input_1150;
      end
      11'b10001111111 : begin
        result = input_1151;
      end
      11'b10010000000 : begin
        result = input_1152;
      end
      11'b10010000001 : begin
        result = input_1153;
      end
      11'b10010000010 : begin
        result = input_1154;
      end
      11'b10010000011 : begin
        result = input_1155;
      end
      11'b10010000100 : begin
        result = input_1156;
      end
      11'b10010000101 : begin
        result = input_1157;
      end
      11'b10010000110 : begin
        result = input_1158;
      end
      11'b10010000111 : begin
        result = input_1159;
      end
      11'b10010001000 : begin
        result = input_1160;
      end
      11'b10010001001 : begin
        result = input_1161;
      end
      11'b10010001010 : begin
        result = input_1162;
      end
      11'b10010001011 : begin
        result = input_1163;
      end
      11'b10010001100 : begin
        result = input_1164;
      end
      11'b10010001101 : begin
        result = input_1165;
      end
      11'b10010001110 : begin
        result = input_1166;
      end
      11'b10010001111 : begin
        result = input_1167;
      end
      11'b10010010000 : begin
        result = input_1168;
      end
      11'b10010010001 : begin
        result = input_1169;
      end
      11'b10010010010 : begin
        result = input_1170;
      end
      11'b10010010011 : begin
        result = input_1171;
      end
      11'b10010010100 : begin
        result = input_1172;
      end
      11'b10010010101 : begin
        result = input_1173;
      end
      11'b10010010110 : begin
        result = input_1174;
      end
      11'b10010010111 : begin
        result = input_1175;
      end
      11'b10010011000 : begin
        result = input_1176;
      end
      11'b10010011001 : begin
        result = input_1177;
      end
      11'b10010011010 : begin
        result = input_1178;
      end
      11'b10010011011 : begin
        result = input_1179;
      end
      11'b10010011100 : begin
        result = input_1180;
      end
      11'b10010011101 : begin
        result = input_1181;
      end
      11'b10010011110 : begin
        result = input_1182;
      end
      11'b10010011111 : begin
        result = input_1183;
      end
      11'b10010100000 : begin
        result = input_1184;
      end
      11'b10010100001 : begin
        result = input_1185;
      end
      11'b10010100010 : begin
        result = input_1186;
      end
      11'b10010100011 : begin
        result = input_1187;
      end
      11'b10010100100 : begin
        result = input_1188;
      end
      11'b10010100101 : begin
        result = input_1189;
      end
      11'b10010100110 : begin
        result = input_1190;
      end
      11'b10010100111 : begin
        result = input_1191;
      end
      11'b10010101000 : begin
        result = input_1192;
      end
      11'b10010101001 : begin
        result = input_1193;
      end
      11'b10010101010 : begin
        result = input_1194;
      end
      11'b10010101011 : begin
        result = input_1195;
      end
      11'b10010101100 : begin
        result = input_1196;
      end
      11'b10010101101 : begin
        result = input_1197;
      end
      11'b10010101110 : begin
        result = input_1198;
      end
      11'b10010101111 : begin
        result = input_1199;
      end
      11'b10010110000 : begin
        result = input_1200;
      end
      11'b10010110001 : begin
        result = input_1201;
      end
      11'b10010110010 : begin
        result = input_1202;
      end
      11'b10010110011 : begin
        result = input_1203;
      end
      11'b10010110100 : begin
        result = input_1204;
      end
      11'b10010110101 : begin
        result = input_1205;
      end
      11'b10010110110 : begin
        result = input_1206;
      end
      11'b10010110111 : begin
        result = input_1207;
      end
      11'b10010111000 : begin
        result = input_1208;
      end
      11'b10010111001 : begin
        result = input_1209;
      end
      11'b10010111010 : begin
        result = input_1210;
      end
      11'b10010111011 : begin
        result = input_1211;
      end
      11'b10010111100 : begin
        result = input_1212;
      end
      11'b10010111101 : begin
        result = input_1213;
      end
      11'b10010111110 : begin
        result = input_1214;
      end
      11'b10010111111 : begin
        result = input_1215;
      end
      11'b10011000000 : begin
        result = input_1216;
      end
      11'b10011000001 : begin
        result = input_1217;
      end
      11'b10011000010 : begin
        result = input_1218;
      end
      11'b10011000011 : begin
        result = input_1219;
      end
      11'b10011000100 : begin
        result = input_1220;
      end
      11'b10011000101 : begin
        result = input_1221;
      end
      11'b10011000110 : begin
        result = input_1222;
      end
      11'b10011000111 : begin
        result = input_1223;
      end
      11'b10011001000 : begin
        result = input_1224;
      end
      11'b10011001001 : begin
        result = input_1225;
      end
      11'b10011001010 : begin
        result = input_1226;
      end
      11'b10011001011 : begin
        result = input_1227;
      end
      11'b10011001100 : begin
        result = input_1228;
      end
      11'b10011001101 : begin
        result = input_1229;
      end
      11'b10011001110 : begin
        result = input_1230;
      end
      11'b10011001111 : begin
        result = input_1231;
      end
      11'b10011010000 : begin
        result = input_1232;
      end
      11'b10011010001 : begin
        result = input_1233;
      end
      11'b10011010010 : begin
        result = input_1234;
      end
      11'b10011010011 : begin
        result = input_1235;
      end
      11'b10011010100 : begin
        result = input_1236;
      end
      11'b10011010101 : begin
        result = input_1237;
      end
      11'b10011010110 : begin
        result = input_1238;
      end
      11'b10011010111 : begin
        result = input_1239;
      end
      11'b10011011000 : begin
        result = input_1240;
      end
      11'b10011011001 : begin
        result = input_1241;
      end
      11'b10011011010 : begin
        result = input_1242;
      end
      11'b10011011011 : begin
        result = input_1243;
      end
      11'b10011011100 : begin
        result = input_1244;
      end
      11'b10011011101 : begin
        result = input_1245;
      end
      11'b10011011110 : begin
        result = input_1246;
      end
      11'b10011011111 : begin
        result = input_1247;
      end
      11'b10011100000 : begin
        result = input_1248;
      end
      11'b10011100001 : begin
        result = input_1249;
      end
      11'b10011100010 : begin
        result = input_1250;
      end
      11'b10011100011 : begin
        result = input_1251;
      end
      11'b10011100100 : begin
        result = input_1252;
      end
      11'b10011100101 : begin
        result = input_1253;
      end
      11'b10011100110 : begin
        result = input_1254;
      end
      11'b10011100111 : begin
        result = input_1255;
      end
      11'b10011101000 : begin
        result = input_1256;
      end
      11'b10011101001 : begin
        result = input_1257;
      end
      11'b10011101010 : begin
        result = input_1258;
      end
      11'b10011101011 : begin
        result = input_1259;
      end
      11'b10011101100 : begin
        result = input_1260;
      end
      11'b10011101101 : begin
        result = input_1261;
      end
      11'b10011101110 : begin
        result = input_1262;
      end
      11'b10011101111 : begin
        result = input_1263;
      end
      11'b10011110000 : begin
        result = input_1264;
      end
      11'b10011110001 : begin
        result = input_1265;
      end
      11'b10011110010 : begin
        result = input_1266;
      end
      11'b10011110011 : begin
        result = input_1267;
      end
      11'b10011110100 : begin
        result = input_1268;
      end
      11'b10011110101 : begin
        result = input_1269;
      end
      11'b10011110110 : begin
        result = input_1270;
      end
      11'b10011110111 : begin
        result = input_1271;
      end
      11'b10011111000 : begin
        result = input_1272;
      end
      11'b10011111001 : begin
        result = input_1273;
      end
      11'b10011111010 : begin
        result = input_1274;
      end
      11'b10011111011 : begin
        result = input_1275;
      end
      11'b10011111100 : begin
        result = input_1276;
      end
      11'b10011111101 : begin
        result = input_1277;
      end
      11'b10011111110 : begin
        result = input_1278;
      end
      11'b10011111111 : begin
        result = input_1279;
      end
      11'b10100000000 : begin
        result = input_1280;
      end
      11'b10100000001 : begin
        result = input_1281;
      end
      11'b10100000010 : begin
        result = input_1282;
      end
      11'b10100000011 : begin
        result = input_1283;
      end
      11'b10100000100 : begin
        result = input_1284;
      end
      11'b10100000101 : begin
        result = input_1285;
      end
      11'b10100000110 : begin
        result = input_1286;
      end
      11'b10100000111 : begin
        result = input_1287;
      end
      11'b10100001000 : begin
        result = input_1288;
      end
      11'b10100001001 : begin
        result = input_1289;
      end
      11'b10100001010 : begin
        result = input_1290;
      end
      11'b10100001011 : begin
        result = input_1291;
      end
      11'b10100001100 : begin
        result = input_1292;
      end
      11'b10100001101 : begin
        result = input_1293;
      end
      11'b10100001110 : begin
        result = input_1294;
      end
      11'b10100001111 : begin
        result = input_1295;
      end
      11'b10100010000 : begin
        result = input_1296;
      end
      11'b10100010001 : begin
        result = input_1297;
      end
      11'b10100010010 : begin
        result = input_1298;
      end
      11'b10100010011 : begin
        result = input_1299;
      end
      11'b10100010100 : begin
        result = input_1300;
      end
      11'b10100010101 : begin
        result = input_1301;
      end
      11'b10100010110 : begin
        result = input_1302;
      end
      11'b10100010111 : begin
        result = input_1303;
      end
      11'b10100011000 : begin
        result = input_1304;
      end
      11'b10100011001 : begin
        result = input_1305;
      end
      11'b10100011010 : begin
        result = input_1306;
      end
      11'b10100011011 : begin
        result = input_1307;
      end
      11'b10100011100 : begin
        result = input_1308;
      end
      11'b10100011101 : begin
        result = input_1309;
      end
      11'b10100011110 : begin
        result = input_1310;
      end
      11'b10100011111 : begin
        result = input_1311;
      end
      11'b10100100000 : begin
        result = input_1312;
      end
      11'b10100100001 : begin
        result = input_1313;
      end
      11'b10100100010 : begin
        result = input_1314;
      end
      11'b10100100011 : begin
        result = input_1315;
      end
      11'b10100100100 : begin
        result = input_1316;
      end
      11'b10100100101 : begin
        result = input_1317;
      end
      11'b10100100110 : begin
        result = input_1318;
      end
      11'b10100100111 : begin
        result = input_1319;
      end
      11'b10100101000 : begin
        result = input_1320;
      end
      11'b10100101001 : begin
        result = input_1321;
      end
      11'b10100101010 : begin
        result = input_1322;
      end
      11'b10100101011 : begin
        result = input_1323;
      end
      11'b10100101100 : begin
        result = input_1324;
      end
      11'b10100101101 : begin
        result = input_1325;
      end
      11'b10100101110 : begin
        result = input_1326;
      end
      11'b10100101111 : begin
        result = input_1327;
      end
      11'b10100110000 : begin
        result = input_1328;
      end
      11'b10100110001 : begin
        result = input_1329;
      end
      11'b10100110010 : begin
        result = input_1330;
      end
      11'b10100110011 : begin
        result = input_1331;
      end
      11'b10100110100 : begin
        result = input_1332;
      end
      11'b10100110101 : begin
        result = input_1333;
      end
      11'b10100110110 : begin
        result = input_1334;
      end
      11'b10100110111 : begin
        result = input_1335;
      end
      11'b10100111000 : begin
        result = input_1336;
      end
      11'b10100111001 : begin
        result = input_1337;
      end
      11'b10100111010 : begin
        result = input_1338;
      end
      11'b10100111011 : begin
        result = input_1339;
      end
      11'b10100111100 : begin
        result = input_1340;
      end
      11'b10100111101 : begin
        result = input_1341;
      end
      11'b10100111110 : begin
        result = input_1342;
      end
      11'b10100111111 : begin
        result = input_1343;
      end
      11'b10101000000 : begin
        result = input_1344;
      end
      11'b10101000001 : begin
        result = input_1345;
      end
      11'b10101000010 : begin
        result = input_1346;
      end
      11'b10101000011 : begin
        result = input_1347;
      end
      11'b10101000100 : begin
        result = input_1348;
      end
      11'b10101000101 : begin
        result = input_1349;
      end
      11'b10101000110 : begin
        result = input_1350;
      end
      11'b10101000111 : begin
        result = input_1351;
      end
      11'b10101001000 : begin
        result = input_1352;
      end
      11'b10101001001 : begin
        result = input_1353;
      end
      11'b10101001010 : begin
        result = input_1354;
      end
      11'b10101001011 : begin
        result = input_1355;
      end
      11'b10101001100 : begin
        result = input_1356;
      end
      11'b10101001101 : begin
        result = input_1357;
      end
      11'b10101001110 : begin
        result = input_1358;
      end
      11'b10101001111 : begin
        result = input_1359;
      end
      11'b10101010000 : begin
        result = input_1360;
      end
      11'b10101010001 : begin
        result = input_1361;
      end
      11'b10101010010 : begin
        result = input_1362;
      end
      11'b10101010011 : begin
        result = input_1363;
      end
      11'b10101010100 : begin
        result = input_1364;
      end
      11'b10101010101 : begin
        result = input_1365;
      end
      11'b10101010110 : begin
        result = input_1366;
      end
      11'b10101010111 : begin
        result = input_1367;
      end
      11'b10101011000 : begin
        result = input_1368;
      end
      11'b10101011001 : begin
        result = input_1369;
      end
      11'b10101011010 : begin
        result = input_1370;
      end
      11'b10101011011 : begin
        result = input_1371;
      end
      11'b10101011100 : begin
        result = input_1372;
      end
      11'b10101011101 : begin
        result = input_1373;
      end
      11'b10101011110 : begin
        result = input_1374;
      end
      11'b10101011111 : begin
        result = input_1375;
      end
      11'b10101100000 : begin
        result = input_1376;
      end
      11'b10101100001 : begin
        result = input_1377;
      end
      11'b10101100010 : begin
        result = input_1378;
      end
      11'b10101100011 : begin
        result = input_1379;
      end
      11'b10101100100 : begin
        result = input_1380;
      end
      11'b10101100101 : begin
        result = input_1381;
      end
      11'b10101100110 : begin
        result = input_1382;
      end
      11'b10101100111 : begin
        result = input_1383;
      end
      11'b10101101000 : begin
        result = input_1384;
      end
      11'b10101101001 : begin
        result = input_1385;
      end
      11'b10101101010 : begin
        result = input_1386;
      end
      11'b10101101011 : begin
        result = input_1387;
      end
      11'b10101101100 : begin
        result = input_1388;
      end
      11'b10101101101 : begin
        result = input_1389;
      end
      11'b10101101110 : begin
        result = input_1390;
      end
      11'b10101101111 : begin
        result = input_1391;
      end
      11'b10101110000 : begin
        result = input_1392;
      end
      11'b10101110001 : begin
        result = input_1393;
      end
      11'b10101110010 : begin
        result = input_1394;
      end
      11'b10101110011 : begin
        result = input_1395;
      end
      11'b10101110100 : begin
        result = input_1396;
      end
      11'b10101110101 : begin
        result = input_1397;
      end
      11'b10101110110 : begin
        result = input_1398;
      end
      11'b10101110111 : begin
        result = input_1399;
      end
      11'b10101111000 : begin
        result = input_1400;
      end
      11'b10101111001 : begin
        result = input_1401;
      end
      11'b10101111010 : begin
        result = input_1402;
      end
      11'b10101111011 : begin
        result = input_1403;
      end
      11'b10101111100 : begin
        result = input_1404;
      end
      11'b10101111101 : begin
        result = input_1405;
      end
      11'b10101111110 : begin
        result = input_1406;
      end
      11'b10101111111 : begin
        result = input_1407;
      end
      11'b10110000000 : begin
        result = input_1408;
      end
      11'b10110000001 : begin
        result = input_1409;
      end
      11'b10110000010 : begin
        result = input_1410;
      end
      11'b10110000011 : begin
        result = input_1411;
      end
      11'b10110000100 : begin
        result = input_1412;
      end
      11'b10110000101 : begin
        result = input_1413;
      end
      11'b10110000110 : begin
        result = input_1414;
      end
      11'b10110000111 : begin
        result = input_1415;
      end
      11'b10110001000 : begin
        result = input_1416;
      end
      11'b10110001001 : begin
        result = input_1417;
      end
      11'b10110001010 : begin
        result = input_1418;
      end
      11'b10110001011 : begin
        result = input_1419;
      end
      11'b10110001100 : begin
        result = input_1420;
      end
      11'b10110001101 : begin
        result = input_1421;
      end
      11'b10110001110 : begin
        result = input_1422;
      end
      11'b10110001111 : begin
        result = input_1423;
      end
      11'b10110010000 : begin
        result = input_1424;
      end
      11'b10110010001 : begin
        result = input_1425;
      end
      11'b10110010010 : begin
        result = input_1426;
      end
      11'b10110010011 : begin
        result = input_1427;
      end
      11'b10110010100 : begin
        result = input_1428;
      end
      11'b10110010101 : begin
        result = input_1429;
      end
      11'b10110010110 : begin
        result = input_1430;
      end
      11'b10110010111 : begin
        result = input_1431;
      end
      11'b10110011000 : begin
        result = input_1432;
      end
      11'b10110011001 : begin
        result = input_1433;
      end
      11'b10110011010 : begin
        result = input_1434;
      end
      11'b10110011011 : begin
        result = input_1435;
      end
      11'b10110011100 : begin
        result = input_1436;
      end
      11'b10110011101 : begin
        result = input_1437;
      end
      11'b10110011110 : begin
        result = input_1438;
      end
      11'b10110011111 : begin
        result = input_1439;
      end
      11'b10110100000 : begin
        result = input_1440;
      end
      11'b10110100001 : begin
        result = input_1441;
      end
      11'b10110100010 : begin
        result = input_1442;
      end
      11'b10110100011 : begin
        result = input_1443;
      end
      11'b10110100100 : begin
        result = input_1444;
      end
      11'b10110100101 : begin
        result = input_1445;
      end
      11'b10110100110 : begin
        result = input_1446;
      end
      11'b10110100111 : begin
        result = input_1447;
      end
      11'b10110101000 : begin
        result = input_1448;
      end
      11'b10110101001 : begin
        result = input_1449;
      end
      11'b10110101010 : begin
        result = input_1450;
      end
      11'b10110101011 : begin
        result = input_1451;
      end
      11'b10110101100 : begin
        result = input_1452;
      end
      11'b10110101101 : begin
        result = input_1453;
      end
      11'b10110101110 : begin
        result = input_1454;
      end
      11'b10110101111 : begin
        result = input_1455;
      end
      11'b10110110000 : begin
        result = input_1456;
      end
      11'b10110110001 : begin
        result = input_1457;
      end
      11'b10110110010 : begin
        result = input_1458;
      end
      11'b10110110011 : begin
        result = input_1459;
      end
      11'b10110110100 : begin
        result = input_1460;
      end
      11'b10110110101 : begin
        result = input_1461;
      end
      11'b10110110110 : begin
        result = input_1462;
      end
      11'b10110110111 : begin
        result = input_1463;
      end
      11'b10110111000 : begin
        result = input_1464;
      end
      11'b10110111001 : begin
        result = input_1465;
      end
      11'b10110111010 : begin
        result = input_1466;
      end
      11'b10110111011 : begin
        result = input_1467;
      end
      11'b10110111100 : begin
        result = input_1468;
      end
      11'b10110111101 : begin
        result = input_1469;
      end
      11'b10110111110 : begin
        result = input_1470;
      end
      11'b10110111111 : begin
        result = input_1471;
      end
      11'b10111000000 : begin
        result = input_1472;
      end
      11'b10111000001 : begin
        result = input_1473;
      end
      11'b10111000010 : begin
        result = input_1474;
      end
      11'b10111000011 : begin
        result = input_1475;
      end
      11'b10111000100 : begin
        result = input_1476;
      end
      11'b10111000101 : begin
        result = input_1477;
      end
      11'b10111000110 : begin
        result = input_1478;
      end
      11'b10111000111 : begin
        result = input_1479;
      end
      11'b10111001000 : begin
        result = input_1480;
      end
      11'b10111001001 : begin
        result = input_1481;
      end
      11'b10111001010 : begin
        result = input_1482;
      end
      11'b10111001011 : begin
        result = input_1483;
      end
      11'b10111001100 : begin
        result = input_1484;
      end
      11'b10111001101 : begin
        result = input_1485;
      end
      11'b10111001110 : begin
        result = input_1486;
      end
      11'b10111001111 : begin
        result = input_1487;
      end
      11'b10111010000 : begin
        result = input_1488;
      end
      11'b10111010001 : begin
        result = input_1489;
      end
      11'b10111010010 : begin
        result = input_1490;
      end
      11'b10111010011 : begin
        result = input_1491;
      end
      11'b10111010100 : begin
        result = input_1492;
      end
      11'b10111010101 : begin
        result = input_1493;
      end
      11'b10111010110 : begin
        result = input_1494;
      end
      11'b10111010111 : begin
        result = input_1495;
      end
      11'b10111011000 : begin
        result = input_1496;
      end
      11'b10111011001 : begin
        result = input_1497;
      end
      11'b10111011010 : begin
        result = input_1498;
      end
      11'b10111011011 : begin
        result = input_1499;
      end
      11'b10111011100 : begin
        result = input_1500;
      end
      11'b10111011101 : begin
        result = input_1501;
      end
      11'b10111011110 : begin
        result = input_1502;
      end
      11'b10111011111 : begin
        result = input_1503;
      end
      11'b10111100000 : begin
        result = input_1504;
      end
      11'b10111100001 : begin
        result = input_1505;
      end
      11'b10111100010 : begin
        result = input_1506;
      end
      11'b10111100011 : begin
        result = input_1507;
      end
      11'b10111100100 : begin
        result = input_1508;
      end
      11'b10111100101 : begin
        result = input_1509;
      end
      11'b10111100110 : begin
        result = input_1510;
      end
      11'b10111100111 : begin
        result = input_1511;
      end
      11'b10111101000 : begin
        result = input_1512;
      end
      11'b10111101001 : begin
        result = input_1513;
      end
      11'b10111101010 : begin
        result = input_1514;
      end
      11'b10111101011 : begin
        result = input_1515;
      end
      11'b10111101100 : begin
        result = input_1516;
      end
      11'b10111101101 : begin
        result = input_1517;
      end
      11'b10111101110 : begin
        result = input_1518;
      end
      11'b10111101111 : begin
        result = input_1519;
      end
      11'b10111110000 : begin
        result = input_1520;
      end
      11'b10111110001 : begin
        result = input_1521;
      end
      11'b10111110010 : begin
        result = input_1522;
      end
      11'b10111110011 : begin
        result = input_1523;
      end
      11'b10111110100 : begin
        result = input_1524;
      end
      11'b10111110101 : begin
        result = input_1525;
      end
      11'b10111110110 : begin
        result = input_1526;
      end
      11'b10111110111 : begin
        result = input_1527;
      end
      11'b10111111000 : begin
        result = input_1528;
      end
      11'b10111111001 : begin
        result = input_1529;
      end
      11'b10111111010 : begin
        result = input_1530;
      end
      11'b10111111011 : begin
        result = input_1531;
      end
      11'b10111111100 : begin
        result = input_1532;
      end
      11'b10111111101 : begin
        result = input_1533;
      end
      11'b10111111110 : begin
        result = input_1534;
      end
      11'b10111111111 : begin
        result = input_1535;
      end
      11'b11000000000 : begin
        result = input_1536;
      end
      11'b11000000001 : begin
        result = input_1537;
      end
      11'b11000000010 : begin
        result = input_1538;
      end
      11'b11000000011 : begin
        result = input_1539;
      end
      11'b11000000100 : begin
        result = input_1540;
      end
      11'b11000000101 : begin
        result = input_1541;
      end
      11'b11000000110 : begin
        result = input_1542;
      end
      11'b11000000111 : begin
        result = input_1543;
      end
      11'b11000001000 : begin
        result = input_1544;
      end
      11'b11000001001 : begin
        result = input_1545;
      end
      11'b11000001010 : begin
        result = input_1546;
      end
      11'b11000001011 : begin
        result = input_1547;
      end
      11'b11000001100 : begin
        result = input_1548;
      end
      11'b11000001101 : begin
        result = input_1549;
      end
      11'b11000001110 : begin
        result = input_1550;
      end
      11'b11000001111 : begin
        result = input_1551;
      end
      11'b11000010000 : begin
        result = input_1552;
      end
      11'b11000010001 : begin
        result = input_1553;
      end
      11'b11000010010 : begin
        result = input_1554;
      end
      11'b11000010011 : begin
        result = input_1555;
      end
      11'b11000010100 : begin
        result = input_1556;
      end
      11'b11000010101 : begin
        result = input_1557;
      end
      11'b11000010110 : begin
        result = input_1558;
      end
      11'b11000010111 : begin
        result = input_1559;
      end
      11'b11000011000 : begin
        result = input_1560;
      end
      11'b11000011001 : begin
        result = input_1561;
      end
      11'b11000011010 : begin
        result = input_1562;
      end
      11'b11000011011 : begin
        result = input_1563;
      end
      11'b11000011100 : begin
        result = input_1564;
      end
      11'b11000011101 : begin
        result = input_1565;
      end
      11'b11000011110 : begin
        result = input_1566;
      end
      11'b11000011111 : begin
        result = input_1567;
      end
      11'b11000100000 : begin
        result = input_1568;
      end
      11'b11000100001 : begin
        result = input_1569;
      end
      11'b11000100010 : begin
        result = input_1570;
      end
      11'b11000100011 : begin
        result = input_1571;
      end
      11'b11000100100 : begin
        result = input_1572;
      end
      11'b11000100101 : begin
        result = input_1573;
      end
      11'b11000100110 : begin
        result = input_1574;
      end
      11'b11000100111 : begin
        result = input_1575;
      end
      11'b11000101000 : begin
        result = input_1576;
      end
      11'b11000101001 : begin
        result = input_1577;
      end
      11'b11000101010 : begin
        result = input_1578;
      end
      11'b11000101011 : begin
        result = input_1579;
      end
      11'b11000101100 : begin
        result = input_1580;
      end
      11'b11000101101 : begin
        result = input_1581;
      end
      11'b11000101110 : begin
        result = input_1582;
      end
      11'b11000101111 : begin
        result = input_1583;
      end
      11'b11000110000 : begin
        result = input_1584;
      end
      11'b11000110001 : begin
        result = input_1585;
      end
      11'b11000110010 : begin
        result = input_1586;
      end
      11'b11000110011 : begin
        result = input_1587;
      end
      11'b11000110100 : begin
        result = input_1588;
      end
      11'b11000110101 : begin
        result = input_1589;
      end
      11'b11000110110 : begin
        result = input_1590;
      end
      11'b11000110111 : begin
        result = input_1591;
      end
      11'b11000111000 : begin
        result = input_1592;
      end
      11'b11000111001 : begin
        result = input_1593;
      end
      11'b11000111010 : begin
        result = input_1594;
      end
      11'b11000111011 : begin
        result = input_1595;
      end
      11'b11000111100 : begin
        result = input_1596;
      end
      11'b11000111101 : begin
        result = input_1597;
      end
      11'b11000111110 : begin
        result = input_1598;
      end
      11'b11000111111 : begin
        result = input_1599;
      end
      11'b11001000000 : begin
        result = input_1600;
      end
      11'b11001000001 : begin
        result = input_1601;
      end
      11'b11001000010 : begin
        result = input_1602;
      end
      11'b11001000011 : begin
        result = input_1603;
      end
      11'b11001000100 : begin
        result = input_1604;
      end
      11'b11001000101 : begin
        result = input_1605;
      end
      11'b11001000110 : begin
        result = input_1606;
      end
      11'b11001000111 : begin
        result = input_1607;
      end
      11'b11001001000 : begin
        result = input_1608;
      end
      11'b11001001001 : begin
        result = input_1609;
      end
      11'b11001001010 : begin
        result = input_1610;
      end
      11'b11001001011 : begin
        result = input_1611;
      end
      11'b11001001100 : begin
        result = input_1612;
      end
      11'b11001001101 : begin
        result = input_1613;
      end
      11'b11001001110 : begin
        result = input_1614;
      end
      11'b11001001111 : begin
        result = input_1615;
      end
      11'b11001010000 : begin
        result = input_1616;
      end
      11'b11001010001 : begin
        result = input_1617;
      end
      11'b11001010010 : begin
        result = input_1618;
      end
      11'b11001010011 : begin
        result = input_1619;
      end
      11'b11001010100 : begin
        result = input_1620;
      end
      11'b11001010101 : begin
        result = input_1621;
      end
      11'b11001010110 : begin
        result = input_1622;
      end
      11'b11001010111 : begin
        result = input_1623;
      end
      11'b11001011000 : begin
        result = input_1624;
      end
      11'b11001011001 : begin
        result = input_1625;
      end
      11'b11001011010 : begin
        result = input_1626;
      end
      11'b11001011011 : begin
        result = input_1627;
      end
      11'b11001011100 : begin
        result = input_1628;
      end
      11'b11001011101 : begin
        result = input_1629;
      end
      11'b11001011110 : begin
        result = input_1630;
      end
      11'b11001011111 : begin
        result = input_1631;
      end
      11'b11001100000 : begin
        result = input_1632;
      end
      11'b11001100001 : begin
        result = input_1633;
      end
      11'b11001100010 : begin
        result = input_1634;
      end
      11'b11001100011 : begin
        result = input_1635;
      end
      11'b11001100100 : begin
        result = input_1636;
      end
      11'b11001100101 : begin
        result = input_1637;
      end
      11'b11001100110 : begin
        result = input_1638;
      end
      11'b11001100111 : begin
        result = input_1639;
      end
      11'b11001101000 : begin
        result = input_1640;
      end
      11'b11001101001 : begin
        result = input_1641;
      end
      11'b11001101010 : begin
        result = input_1642;
      end
      11'b11001101011 : begin
        result = input_1643;
      end
      11'b11001101100 : begin
        result = input_1644;
      end
      11'b11001101101 : begin
        result = input_1645;
      end
      11'b11001101110 : begin
        result = input_1646;
      end
      11'b11001101111 : begin
        result = input_1647;
      end
      11'b11001110000 : begin
        result = input_1648;
      end
      11'b11001110001 : begin
        result = input_1649;
      end
      11'b11001110010 : begin
        result = input_1650;
      end
      11'b11001110011 : begin
        result = input_1651;
      end
      11'b11001110100 : begin
        result = input_1652;
      end
      11'b11001110101 : begin
        result = input_1653;
      end
      11'b11001110110 : begin
        result = input_1654;
      end
      11'b11001110111 : begin
        result = input_1655;
      end
      11'b11001111000 : begin
        result = input_1656;
      end
      11'b11001111001 : begin
        result = input_1657;
      end
      11'b11001111010 : begin
        result = input_1658;
      end
      11'b11001111011 : begin
        result = input_1659;
      end
      11'b11001111100 : begin
        result = input_1660;
      end
      11'b11001111101 : begin
        result = input_1661;
      end
      11'b11001111110 : begin
        result = input_1662;
      end
      11'b11001111111 : begin
        result = input_1663;
      end
      11'b11010000000 : begin
        result = input_1664;
      end
      11'b11010000001 : begin
        result = input_1665;
      end
      11'b11010000010 : begin
        result = input_1666;
      end
      11'b11010000011 : begin
        result = input_1667;
      end
      11'b11010000100 : begin
        result = input_1668;
      end
      11'b11010000101 : begin
        result = input_1669;
      end
      11'b11010000110 : begin
        result = input_1670;
      end
      11'b11010000111 : begin
        result = input_1671;
      end
      11'b11010001000 : begin
        result = input_1672;
      end
      11'b11010001001 : begin
        result = input_1673;
      end
      11'b11010001010 : begin
        result = input_1674;
      end
      11'b11010001011 : begin
        result = input_1675;
      end
      11'b11010001100 : begin
        result = input_1676;
      end
      11'b11010001101 : begin
        result = input_1677;
      end
      11'b11010001110 : begin
        result = input_1678;
      end
      11'b11010001111 : begin
        result = input_1679;
      end
      11'b11010010000 : begin
        result = input_1680;
      end
      11'b11010010001 : begin
        result = input_1681;
      end
      11'b11010010010 : begin
        result = input_1682;
      end
      11'b11010010011 : begin
        result = input_1683;
      end
      11'b11010010100 : begin
        result = input_1684;
      end
      11'b11010010101 : begin
        result = input_1685;
      end
      11'b11010010110 : begin
        result = input_1686;
      end
      11'b11010010111 : begin
        result = input_1687;
      end
      11'b11010011000 : begin
        result = input_1688;
      end
      11'b11010011001 : begin
        result = input_1689;
      end
      11'b11010011010 : begin
        result = input_1690;
      end
      11'b11010011011 : begin
        result = input_1691;
      end
      11'b11010011100 : begin
        result = input_1692;
      end
      11'b11010011101 : begin
        result = input_1693;
      end
      11'b11010011110 : begin
        result = input_1694;
      end
      11'b11010011111 : begin
        result = input_1695;
      end
      11'b11010100000 : begin
        result = input_1696;
      end
      11'b11010100001 : begin
        result = input_1697;
      end
      11'b11010100010 : begin
        result = input_1698;
      end
      11'b11010100011 : begin
        result = input_1699;
      end
      11'b11010100100 : begin
        result = input_1700;
      end
      11'b11010100101 : begin
        result = input_1701;
      end
      11'b11010100110 : begin
        result = input_1702;
      end
      11'b11010100111 : begin
        result = input_1703;
      end
      11'b11010101000 : begin
        result = input_1704;
      end
      11'b11010101001 : begin
        result = input_1705;
      end
      11'b11010101010 : begin
        result = input_1706;
      end
      11'b11010101011 : begin
        result = input_1707;
      end
      11'b11010101100 : begin
        result = input_1708;
      end
      11'b11010101101 : begin
        result = input_1709;
      end
      11'b11010101110 : begin
        result = input_1710;
      end
      11'b11010101111 : begin
        result = input_1711;
      end
      11'b11010110000 : begin
        result = input_1712;
      end
      11'b11010110001 : begin
        result = input_1713;
      end
      11'b11010110010 : begin
        result = input_1714;
      end
      11'b11010110011 : begin
        result = input_1715;
      end
      11'b11010110100 : begin
        result = input_1716;
      end
      11'b11010110101 : begin
        result = input_1717;
      end
      11'b11010110110 : begin
        result = input_1718;
      end
      11'b11010110111 : begin
        result = input_1719;
      end
      11'b11010111000 : begin
        result = input_1720;
      end
      11'b11010111001 : begin
        result = input_1721;
      end
      11'b11010111010 : begin
        result = input_1722;
      end
      11'b11010111011 : begin
        result = input_1723;
      end
      11'b11010111100 : begin
        result = input_1724;
      end
      11'b11010111101 : begin
        result = input_1725;
      end
      11'b11010111110 : begin
        result = input_1726;
      end
      11'b11010111111 : begin
        result = input_1727;
      end
      11'b11011000000 : begin
        result = input_1728;
      end
      11'b11011000001 : begin
        result = input_1729;
      end
      11'b11011000010 : begin
        result = input_1730;
      end
      11'b11011000011 : begin
        result = input_1731;
      end
      11'b11011000100 : begin
        result = input_1732;
      end
      11'b11011000101 : begin
        result = input_1733;
      end
      11'b11011000110 : begin
        result = input_1734;
      end
      11'b11011000111 : begin
        result = input_1735;
      end
      11'b11011001000 : begin
        result = input_1736;
      end
      11'b11011001001 : begin
        result = input_1737;
      end
      11'b11011001010 : begin
        result = input_1738;
      end
      11'b11011001011 : begin
        result = input_1739;
      end
      11'b11011001100 : begin
        result = input_1740;
      end
      11'b11011001101 : begin
        result = input_1741;
      end
      11'b11011001110 : begin
        result = input_1742;
      end
      11'b11011001111 : begin
        result = input_1743;
      end
      11'b11011010000 : begin
        result = input_1744;
      end
      11'b11011010001 : begin
        result = input_1745;
      end
      11'b11011010010 : begin
        result = input_1746;
      end
      11'b11011010011 : begin
        result = input_1747;
      end
      11'b11011010100 : begin
        result = input_1748;
      end
      11'b11011010101 : begin
        result = input_1749;
      end
      11'b11011010110 : begin
        result = input_1750;
      end
      11'b11011010111 : begin
        result = input_1751;
      end
      11'b11011011000 : begin
        result = input_1752;
      end
      11'b11011011001 : begin
        result = input_1753;
      end
      11'b11011011010 : begin
        result = input_1754;
      end
      11'b11011011011 : begin
        result = input_1755;
      end
      11'b11011011100 : begin
        result = input_1756;
      end
      11'b11011011101 : begin
        result = input_1757;
      end
      11'b11011011110 : begin
        result = input_1758;
      end
      11'b11011011111 : begin
        result = input_1759;
      end
      11'b11011100000 : begin
        result = input_1760;
      end
      11'b11011100001 : begin
        result = input_1761;
      end
      11'b11011100010 : begin
        result = input_1762;
      end
      11'b11011100011 : begin
        result = input_1763;
      end
      11'b11011100100 : begin
        result = input_1764;
      end
      11'b11011100101 : begin
        result = input_1765;
      end
      11'b11011100110 : begin
        result = input_1766;
      end
      11'b11011100111 : begin
        result = input_1767;
      end
      11'b11011101000 : begin
        result = input_1768;
      end
      11'b11011101001 : begin
        result = input_1769;
      end
      11'b11011101010 : begin
        result = input_1770;
      end
      11'b11011101011 : begin
        result = input_1771;
      end
      11'b11011101100 : begin
        result = input_1772;
      end
      11'b11011101101 : begin
        result = input_1773;
      end
      11'b11011101110 : begin
        result = input_1774;
      end
      11'b11011101111 : begin
        result = input_1775;
      end
      11'b11011110000 : begin
        result = input_1776;
      end
      11'b11011110001 : begin
        result = input_1777;
      end
      11'b11011110010 : begin
        result = input_1778;
      end
      11'b11011110011 : begin
        result = input_1779;
      end
      11'b11011110100 : begin
        result = input_1780;
      end
      11'b11011110101 : begin
        result = input_1781;
      end
      11'b11011110110 : begin
        result = input_1782;
      end
      11'b11011110111 : begin
        result = input_1783;
      end
      11'b11011111000 : begin
        result = input_1784;
      end
      11'b11011111001 : begin
        result = input_1785;
      end
      11'b11011111010 : begin
        result = input_1786;
      end
      11'b11011111011 : begin
        result = input_1787;
      end
      11'b11011111100 : begin
        result = input_1788;
      end
      11'b11011111101 : begin
        result = input_1789;
      end
      11'b11011111110 : begin
        result = input_1790;
      end
      11'b11011111111 : begin
        result = input_1791;
      end
      11'b11100000000 : begin
        result = input_1792;
      end
      11'b11100000001 : begin
        result = input_1793;
      end
      11'b11100000010 : begin
        result = input_1794;
      end
      11'b11100000011 : begin
        result = input_1795;
      end
      11'b11100000100 : begin
        result = input_1796;
      end
      11'b11100000101 : begin
        result = input_1797;
      end
      11'b11100000110 : begin
        result = input_1798;
      end
      11'b11100000111 : begin
        result = input_1799;
      end
      11'b11100001000 : begin
        result = input_1800;
      end
      11'b11100001001 : begin
        result = input_1801;
      end
      11'b11100001010 : begin
        result = input_1802;
      end
      11'b11100001011 : begin
        result = input_1803;
      end
      11'b11100001100 : begin
        result = input_1804;
      end
      11'b11100001101 : begin
        result = input_1805;
      end
      11'b11100001110 : begin
        result = input_1806;
      end
      11'b11100001111 : begin
        result = input_1807;
      end
      11'b11100010000 : begin
        result = input_1808;
      end
      11'b11100010001 : begin
        result = input_1809;
      end
      11'b11100010010 : begin
        result = input_1810;
      end
      11'b11100010011 : begin
        result = input_1811;
      end
      11'b11100010100 : begin
        result = input_1812;
      end
      11'b11100010101 : begin
        result = input_1813;
      end
      11'b11100010110 : begin
        result = input_1814;
      end
      11'b11100010111 : begin
        result = input_1815;
      end
      11'b11100011000 : begin
        result = input_1816;
      end
      11'b11100011001 : begin
        result = input_1817;
      end
      11'b11100011010 : begin
        result = input_1818;
      end
      11'b11100011011 : begin
        result = input_1819;
      end
      11'b11100011100 : begin
        result = input_1820;
      end
      11'b11100011101 : begin
        result = input_1821;
      end
      11'b11100011110 : begin
        result = input_1822;
      end
      11'b11100011111 : begin
        result = input_1823;
      end
      11'b11100100000 : begin
        result = input_1824;
      end
      11'b11100100001 : begin
        result = input_1825;
      end
      11'b11100100010 : begin
        result = input_1826;
      end
      11'b11100100011 : begin
        result = input_1827;
      end
      11'b11100100100 : begin
        result = input_1828;
      end
      11'b11100100101 : begin
        result = input_1829;
      end
      11'b11100100110 : begin
        result = input_1830;
      end
      11'b11100100111 : begin
        result = input_1831;
      end
      11'b11100101000 : begin
        result = input_1832;
      end
      11'b11100101001 : begin
        result = input_1833;
      end
      11'b11100101010 : begin
        result = input_1834;
      end
      11'b11100101011 : begin
        result = input_1835;
      end
      11'b11100101100 : begin
        result = input_1836;
      end
      11'b11100101101 : begin
        result = input_1837;
      end
      11'b11100101110 : begin
        result = input_1838;
      end
      11'b11100101111 : begin
        result = input_1839;
      end
      11'b11100110000 : begin
        result = input_1840;
      end
      11'b11100110001 : begin
        result = input_1841;
      end
      11'b11100110010 : begin
        result = input_1842;
      end
      11'b11100110011 : begin
        result = input_1843;
      end
      11'b11100110100 : begin
        result = input_1844;
      end
      11'b11100110101 : begin
        result = input_1845;
      end
      11'b11100110110 : begin
        result = input_1846;
      end
      11'b11100110111 : begin
        result = input_1847;
      end
      11'b11100111000 : begin
        result = input_1848;
      end
      11'b11100111001 : begin
        result = input_1849;
      end
      11'b11100111010 : begin
        result = input_1850;
      end
      11'b11100111011 : begin
        result = input_1851;
      end
      11'b11100111100 : begin
        result = input_1852;
      end
      11'b11100111101 : begin
        result = input_1853;
      end
      11'b11100111110 : begin
        result = input_1854;
      end
      11'b11100111111 : begin
        result = input_1855;
      end
      11'b11101000000 : begin
        result = input_1856;
      end
      11'b11101000001 : begin
        result = input_1857;
      end
      11'b11101000010 : begin
        result = input_1858;
      end
      11'b11101000011 : begin
        result = input_1859;
      end
      11'b11101000100 : begin
        result = input_1860;
      end
      11'b11101000101 : begin
        result = input_1861;
      end
      11'b11101000110 : begin
        result = input_1862;
      end
      11'b11101000111 : begin
        result = input_1863;
      end
      11'b11101001000 : begin
        result = input_1864;
      end
      11'b11101001001 : begin
        result = input_1865;
      end
      11'b11101001010 : begin
        result = input_1866;
      end
      11'b11101001011 : begin
        result = input_1867;
      end
      11'b11101001100 : begin
        result = input_1868;
      end
      11'b11101001101 : begin
        result = input_1869;
      end
      11'b11101001110 : begin
        result = input_1870;
      end
      11'b11101001111 : begin
        result = input_1871;
      end
      11'b11101010000 : begin
        result = input_1872;
      end
      11'b11101010001 : begin
        result = input_1873;
      end
      11'b11101010010 : begin
        result = input_1874;
      end
      11'b11101010011 : begin
        result = input_1875;
      end
      11'b11101010100 : begin
        result = input_1876;
      end
      11'b11101010101 : begin
        result = input_1877;
      end
      11'b11101010110 : begin
        result = input_1878;
      end
      11'b11101010111 : begin
        result = input_1879;
      end
      11'b11101011000 : begin
        result = input_1880;
      end
      11'b11101011001 : begin
        result = input_1881;
      end
      11'b11101011010 : begin
        result = input_1882;
      end
      11'b11101011011 : begin
        result = input_1883;
      end
      11'b11101011100 : begin
        result = input_1884;
      end
      11'b11101011101 : begin
        result = input_1885;
      end
      11'b11101011110 : begin
        result = input_1886;
      end
      11'b11101011111 : begin
        result = input_1887;
      end
      11'b11101100000 : begin
        result = input_1888;
      end
      11'b11101100001 : begin
        result = input_1889;
      end
      11'b11101100010 : begin
        result = input_1890;
      end
      11'b11101100011 : begin
        result = input_1891;
      end
      11'b11101100100 : begin
        result = input_1892;
      end
      11'b11101100101 : begin
        result = input_1893;
      end
      11'b11101100110 : begin
        result = input_1894;
      end
      11'b11101100111 : begin
        result = input_1895;
      end
      11'b11101101000 : begin
        result = input_1896;
      end
      11'b11101101001 : begin
        result = input_1897;
      end
      11'b11101101010 : begin
        result = input_1898;
      end
      11'b11101101011 : begin
        result = input_1899;
      end
      11'b11101101100 : begin
        result = input_1900;
      end
      11'b11101101101 : begin
        result = input_1901;
      end
      11'b11101101110 : begin
        result = input_1902;
      end
      11'b11101101111 : begin
        result = input_1903;
      end
      11'b11101110000 : begin
        result = input_1904;
      end
      11'b11101110001 : begin
        result = input_1905;
      end
      11'b11101110010 : begin
        result = input_1906;
      end
      11'b11101110011 : begin
        result = input_1907;
      end
      11'b11101110100 : begin
        result = input_1908;
      end
      11'b11101110101 : begin
        result = input_1909;
      end
      11'b11101110110 : begin
        result = input_1910;
      end
      11'b11101110111 : begin
        result = input_1911;
      end
      11'b11101111000 : begin
        result = input_1912;
      end
      11'b11101111001 : begin
        result = input_1913;
      end
      11'b11101111010 : begin
        result = input_1914;
      end
      11'b11101111011 : begin
        result = input_1915;
      end
      11'b11101111100 : begin
        result = input_1916;
      end
      11'b11101111101 : begin
        result = input_1917;
      end
      11'b11101111110 : begin
        result = input_1918;
      end
      11'b11101111111 : begin
        result = input_1919;
      end
      11'b11110000000 : begin
        result = input_1920;
      end
      11'b11110000001 : begin
        result = input_1921;
      end
      11'b11110000010 : begin
        result = input_1922;
      end
      11'b11110000011 : begin
        result = input_1923;
      end
      11'b11110000100 : begin
        result = input_1924;
      end
      11'b11110000101 : begin
        result = input_1925;
      end
      11'b11110000110 : begin
        result = input_1926;
      end
      11'b11110000111 : begin
        result = input_1927;
      end
      11'b11110001000 : begin
        result = input_1928;
      end
      11'b11110001001 : begin
        result = input_1929;
      end
      11'b11110001010 : begin
        result = input_1930;
      end
      11'b11110001011 : begin
        result = input_1931;
      end
      11'b11110001100 : begin
        result = input_1932;
      end
      11'b11110001101 : begin
        result = input_1933;
      end
      11'b11110001110 : begin
        result = input_1934;
      end
      11'b11110001111 : begin
        result = input_1935;
      end
      11'b11110010000 : begin
        result = input_1936;
      end
      11'b11110010001 : begin
        result = input_1937;
      end
      11'b11110010010 : begin
        result = input_1938;
      end
      11'b11110010011 : begin
        result = input_1939;
      end
      11'b11110010100 : begin
        result = input_1940;
      end
      11'b11110010101 : begin
        result = input_1941;
      end
      11'b11110010110 : begin
        result = input_1942;
      end
      11'b11110010111 : begin
        result = input_1943;
      end
      11'b11110011000 : begin
        result = input_1944;
      end
      11'b11110011001 : begin
        result = input_1945;
      end
      11'b11110011010 : begin
        result = input_1946;
      end
      11'b11110011011 : begin
        result = input_1947;
      end
      11'b11110011100 : begin
        result = input_1948;
      end
      11'b11110011101 : begin
        result = input_1949;
      end
      11'b11110011110 : begin
        result = input_1950;
      end
      11'b11110011111 : begin
        result = input_1951;
      end
      11'b11110100000 : begin
        result = input_1952;
      end
      11'b11110100001 : begin
        result = input_1953;
      end
      11'b11110100010 : begin
        result = input_1954;
      end
      11'b11110100011 : begin
        result = input_1955;
      end
      11'b11110100100 : begin
        result = input_1956;
      end
      11'b11110100101 : begin
        result = input_1957;
      end
      11'b11110100110 : begin
        result = input_1958;
      end
      11'b11110100111 : begin
        result = input_1959;
      end
      11'b11110101000 : begin
        result = input_1960;
      end
      11'b11110101001 : begin
        result = input_1961;
      end
      11'b11110101010 : begin
        result = input_1962;
      end
      11'b11110101011 : begin
        result = input_1963;
      end
      11'b11110101100 : begin
        result = input_1964;
      end
      11'b11110101101 : begin
        result = input_1965;
      end
      11'b11110101110 : begin
        result = input_1966;
      end
      11'b11110101111 : begin
        result = input_1967;
      end
      11'b11110110000 : begin
        result = input_1968;
      end
      11'b11110110001 : begin
        result = input_1969;
      end
      11'b11110110010 : begin
        result = input_1970;
      end
      11'b11110110011 : begin
        result = input_1971;
      end
      11'b11110110100 : begin
        result = input_1972;
      end
      11'b11110110101 : begin
        result = input_1973;
      end
      11'b11110110110 : begin
        result = input_1974;
      end
      11'b11110110111 : begin
        result = input_1975;
      end
      11'b11110111000 : begin
        result = input_1976;
      end
      11'b11110111001 : begin
        result = input_1977;
      end
      11'b11110111010 : begin
        result = input_1978;
      end
      11'b11110111011 : begin
        result = input_1979;
      end
      11'b11110111100 : begin
        result = input_1980;
      end
      11'b11110111101 : begin
        result = input_1981;
      end
      11'b11110111110 : begin
        result = input_1982;
      end
      11'b11110111111 : begin
        result = input_1983;
      end
      11'b11111000000 : begin
        result = input_1984;
      end
      11'b11111000001 : begin
        result = input_1985;
      end
      11'b11111000010 : begin
        result = input_1986;
      end
      11'b11111000011 : begin
        result = input_1987;
      end
      11'b11111000100 : begin
        result = input_1988;
      end
      11'b11111000101 : begin
        result = input_1989;
      end
      11'b11111000110 : begin
        result = input_1990;
      end
      11'b11111000111 : begin
        result = input_1991;
      end
      11'b11111001000 : begin
        result = input_1992;
      end
      11'b11111001001 : begin
        result = input_1993;
      end
      11'b11111001010 : begin
        result = input_1994;
      end
      11'b11111001011 : begin
        result = input_1995;
      end
      11'b11111001100 : begin
        result = input_1996;
      end
      11'b11111001101 : begin
        result = input_1997;
      end
      11'b11111001110 : begin
        result = input_1998;
      end
      11'b11111001111 : begin
        result = input_1999;
      end
      11'b11111010000 : begin
        result = input_2000;
      end
      11'b11111010001 : begin
        result = input_2001;
      end
      11'b11111010010 : begin
        result = input_2002;
      end
      11'b11111010011 : begin
        result = input_2003;
      end
      11'b11111010100 : begin
        result = input_2004;
      end
      11'b11111010101 : begin
        result = input_2005;
      end
      11'b11111010110 : begin
        result = input_2006;
      end
      11'b11111010111 : begin
        result = input_2007;
      end
      11'b11111011000 : begin
        result = input_2008;
      end
      11'b11111011001 : begin
        result = input_2009;
      end
      11'b11111011010 : begin
        result = input_2010;
      end
      11'b11111011011 : begin
        result = input_2011;
      end
      11'b11111011100 : begin
        result = input_2012;
      end
      11'b11111011101 : begin
        result = input_2013;
      end
      11'b11111011110 : begin
        result = input_2014;
      end
      11'b11111011111 : begin
        result = input_2015;
      end
      11'b11111100000 : begin
        result = input_2016;
      end
      11'b11111100001 : begin
        result = input_2017;
      end
      11'b11111100010 : begin
        result = input_2018;
      end
      11'b11111100011 : begin
        result = input_2019;
      end
      11'b11111100100 : begin
        result = input_2020;
      end
      11'b11111100101 : begin
        result = input_2021;
      end
      11'b11111100110 : begin
        result = input_2022;
      end
      11'b11111100111 : begin
        result = input_2023;
      end
      11'b11111101000 : begin
        result = input_2024;
      end
      11'b11111101001 : begin
        result = input_2025;
      end
      11'b11111101010 : begin
        result = input_2026;
      end
      11'b11111101011 : begin
        result = input_2027;
      end
      11'b11111101100 : begin
        result = input_2028;
      end
      11'b11111101101 : begin
        result = input_2029;
      end
      11'b11111101110 : begin
        result = input_2030;
      end
      11'b11111101111 : begin
        result = input_2031;
      end
      11'b11111110000 : begin
        result = input_2032;
      end
      11'b11111110001 : begin
        result = input_2033;
      end
      11'b11111110010 : begin
        result = input_2034;
      end
      11'b11111110011 : begin
        result = input_2035;
      end
      11'b11111110100 : begin
        result = input_2036;
      end
      11'b11111110101 : begin
        result = input_2037;
      end
      11'b11111110110 : begin
        result = input_2038;
      end
      11'b11111110111 : begin
        result = input_2039;
      end
      11'b11111111000 : begin
        result = input_2040;
      end
      11'b11111111001 : begin
        result = input_2041;
      end
      11'b11111111010 : begin
        result = input_2042;
      end
      11'b11111111011 : begin
        result = input_2043;
      end
      11'b11111111100 : begin
        result = input_2044;
      end
      11'b11111111101 : begin
        result = input_2045;
      end
      11'b11111111110 : begin
        result = input_2046;
      end
      default : begin
        result = input_2047;
      end
    endcase
    MUX_v_5_2048_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i9_1o3_0cffcd7ae8128c5cac71e8022405e1ebb1_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Sat Nov  2 10:26:21 2019
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i9_1o3_0cffcd7ae8128c5cac71e8022405e1ebb1
// ------------------------------------------------------------------


module ROM_1i9_1o3_0cffcd7ae8128c5cac71e8022405e1ebb1 (
  I_1, O_1
);
  input [8:0] I_1;
  output [2:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_3_320_2(3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000,
      3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000,
      3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000,
      3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000,
      3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000,
      3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000,
      3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001,
      3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001,
      3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001,
      3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001,
      3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001,
      3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001,
      3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001,
      3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010,
      3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010,
      3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010,
      3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010,
      3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010,
      3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010,
      3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011,
      3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011,
      3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011,
      3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011,
      3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011,
      3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011,
      3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b100,
      3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
      3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
      3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
      3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
      3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
      3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
      3'b100, 3'b100, 3'b100, I_1);

  function automatic [2:0] MUX_v_3_320_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [2:0] input_2;
    input [2:0] input_3;
    input [2:0] input_4;
    input [2:0] input_5;
    input [2:0] input_6;
    input [2:0] input_7;
    input [2:0] input_8;
    input [2:0] input_9;
    input [2:0] input_10;
    input [2:0] input_11;
    input [2:0] input_12;
    input [2:0] input_13;
    input [2:0] input_14;
    input [2:0] input_15;
    input [2:0] input_16;
    input [2:0] input_17;
    input [2:0] input_18;
    input [2:0] input_19;
    input [2:0] input_20;
    input [2:0] input_21;
    input [2:0] input_22;
    input [2:0] input_23;
    input [2:0] input_24;
    input [2:0] input_25;
    input [2:0] input_26;
    input [2:0] input_27;
    input [2:0] input_28;
    input [2:0] input_29;
    input [2:0] input_30;
    input [2:0] input_31;
    input [2:0] input_32;
    input [2:0] input_33;
    input [2:0] input_34;
    input [2:0] input_35;
    input [2:0] input_36;
    input [2:0] input_37;
    input [2:0] input_38;
    input [2:0] input_39;
    input [2:0] input_40;
    input [2:0] input_41;
    input [2:0] input_42;
    input [2:0] input_43;
    input [2:0] input_44;
    input [2:0] input_45;
    input [2:0] input_46;
    input [2:0] input_47;
    input [2:0] input_48;
    input [2:0] input_49;
    input [2:0] input_50;
    input [2:0] input_51;
    input [2:0] input_52;
    input [2:0] input_53;
    input [2:0] input_54;
    input [2:0] input_55;
    input [2:0] input_56;
    input [2:0] input_57;
    input [2:0] input_58;
    input [2:0] input_59;
    input [2:0] input_60;
    input [2:0] input_61;
    input [2:0] input_62;
    input [2:0] input_63;
    input [2:0] input_64;
    input [2:0] input_65;
    input [2:0] input_66;
    input [2:0] input_67;
    input [2:0] input_68;
    input [2:0] input_69;
    input [2:0] input_70;
    input [2:0] input_71;
    input [2:0] input_72;
    input [2:0] input_73;
    input [2:0] input_74;
    input [2:0] input_75;
    input [2:0] input_76;
    input [2:0] input_77;
    input [2:0] input_78;
    input [2:0] input_79;
    input [2:0] input_80;
    input [2:0] input_81;
    input [2:0] input_82;
    input [2:0] input_83;
    input [2:0] input_84;
    input [2:0] input_85;
    input [2:0] input_86;
    input [2:0] input_87;
    input [2:0] input_88;
    input [2:0] input_89;
    input [2:0] input_90;
    input [2:0] input_91;
    input [2:0] input_92;
    input [2:0] input_93;
    input [2:0] input_94;
    input [2:0] input_95;
    input [2:0] input_96;
    input [2:0] input_97;
    input [2:0] input_98;
    input [2:0] input_99;
    input [2:0] input_100;
    input [2:0] input_101;
    input [2:0] input_102;
    input [2:0] input_103;
    input [2:0] input_104;
    input [2:0] input_105;
    input [2:0] input_106;
    input [2:0] input_107;
    input [2:0] input_108;
    input [2:0] input_109;
    input [2:0] input_110;
    input [2:0] input_111;
    input [2:0] input_112;
    input [2:0] input_113;
    input [2:0] input_114;
    input [2:0] input_115;
    input [2:0] input_116;
    input [2:0] input_117;
    input [2:0] input_118;
    input [2:0] input_119;
    input [2:0] input_120;
    input [2:0] input_121;
    input [2:0] input_122;
    input [2:0] input_123;
    input [2:0] input_124;
    input [2:0] input_125;
    input [2:0] input_126;
    input [2:0] input_127;
    input [2:0] input_128;
    input [2:0] input_129;
    input [2:0] input_130;
    input [2:0] input_131;
    input [2:0] input_132;
    input [2:0] input_133;
    input [2:0] input_134;
    input [2:0] input_135;
    input [2:0] input_136;
    input [2:0] input_137;
    input [2:0] input_138;
    input [2:0] input_139;
    input [2:0] input_140;
    input [2:0] input_141;
    input [2:0] input_142;
    input [2:0] input_143;
    input [2:0] input_144;
    input [2:0] input_145;
    input [2:0] input_146;
    input [2:0] input_147;
    input [2:0] input_148;
    input [2:0] input_149;
    input [2:0] input_150;
    input [2:0] input_151;
    input [2:0] input_152;
    input [2:0] input_153;
    input [2:0] input_154;
    input [2:0] input_155;
    input [2:0] input_156;
    input [2:0] input_157;
    input [2:0] input_158;
    input [2:0] input_159;
    input [2:0] input_160;
    input [2:0] input_161;
    input [2:0] input_162;
    input [2:0] input_163;
    input [2:0] input_164;
    input [2:0] input_165;
    input [2:0] input_166;
    input [2:0] input_167;
    input [2:0] input_168;
    input [2:0] input_169;
    input [2:0] input_170;
    input [2:0] input_171;
    input [2:0] input_172;
    input [2:0] input_173;
    input [2:0] input_174;
    input [2:0] input_175;
    input [2:0] input_176;
    input [2:0] input_177;
    input [2:0] input_178;
    input [2:0] input_179;
    input [2:0] input_180;
    input [2:0] input_181;
    input [2:0] input_182;
    input [2:0] input_183;
    input [2:0] input_184;
    input [2:0] input_185;
    input [2:0] input_186;
    input [2:0] input_187;
    input [2:0] input_188;
    input [2:0] input_189;
    input [2:0] input_190;
    input [2:0] input_191;
    input [2:0] input_192;
    input [2:0] input_193;
    input [2:0] input_194;
    input [2:0] input_195;
    input [2:0] input_196;
    input [2:0] input_197;
    input [2:0] input_198;
    input [2:0] input_199;
    input [2:0] input_200;
    input [2:0] input_201;
    input [2:0] input_202;
    input [2:0] input_203;
    input [2:0] input_204;
    input [2:0] input_205;
    input [2:0] input_206;
    input [2:0] input_207;
    input [2:0] input_208;
    input [2:0] input_209;
    input [2:0] input_210;
    input [2:0] input_211;
    input [2:0] input_212;
    input [2:0] input_213;
    input [2:0] input_214;
    input [2:0] input_215;
    input [2:0] input_216;
    input [2:0] input_217;
    input [2:0] input_218;
    input [2:0] input_219;
    input [2:0] input_220;
    input [2:0] input_221;
    input [2:0] input_222;
    input [2:0] input_223;
    input [2:0] input_224;
    input [2:0] input_225;
    input [2:0] input_226;
    input [2:0] input_227;
    input [2:0] input_228;
    input [2:0] input_229;
    input [2:0] input_230;
    input [2:0] input_231;
    input [2:0] input_232;
    input [2:0] input_233;
    input [2:0] input_234;
    input [2:0] input_235;
    input [2:0] input_236;
    input [2:0] input_237;
    input [2:0] input_238;
    input [2:0] input_239;
    input [2:0] input_240;
    input [2:0] input_241;
    input [2:0] input_242;
    input [2:0] input_243;
    input [2:0] input_244;
    input [2:0] input_245;
    input [2:0] input_246;
    input [2:0] input_247;
    input [2:0] input_248;
    input [2:0] input_249;
    input [2:0] input_250;
    input [2:0] input_251;
    input [2:0] input_252;
    input [2:0] input_253;
    input [2:0] input_254;
    input [2:0] input_255;
    input [2:0] input_256;
    input [2:0] input_257;
    input [2:0] input_258;
    input [2:0] input_259;
    input [2:0] input_260;
    input [2:0] input_261;
    input [2:0] input_262;
    input [2:0] input_263;
    input [2:0] input_264;
    input [2:0] input_265;
    input [2:0] input_266;
    input [2:0] input_267;
    input [2:0] input_268;
    input [2:0] input_269;
    input [2:0] input_270;
    input [2:0] input_271;
    input [2:0] input_272;
    input [2:0] input_273;
    input [2:0] input_274;
    input [2:0] input_275;
    input [2:0] input_276;
    input [2:0] input_277;
    input [2:0] input_278;
    input [2:0] input_279;
    input [2:0] input_280;
    input [2:0] input_281;
    input [2:0] input_282;
    input [2:0] input_283;
    input [2:0] input_284;
    input [2:0] input_285;
    input [2:0] input_286;
    input [2:0] input_287;
    input [2:0] input_288;
    input [2:0] input_289;
    input [2:0] input_290;
    input [2:0] input_291;
    input [2:0] input_292;
    input [2:0] input_293;
    input [2:0] input_294;
    input [2:0] input_295;
    input [2:0] input_296;
    input [2:0] input_297;
    input [2:0] input_298;
    input [2:0] input_299;
    input [2:0] input_300;
    input [2:0] input_301;
    input [2:0] input_302;
    input [2:0] input_303;
    input [2:0] input_304;
    input [2:0] input_305;
    input [2:0] input_306;
    input [2:0] input_307;
    input [2:0] input_308;
    input [2:0] input_309;
    input [2:0] input_310;
    input [2:0] input_311;
    input [2:0] input_312;
    input [2:0] input_313;
    input [2:0] input_314;
    input [2:0] input_315;
    input [2:0] input_316;
    input [2:0] input_317;
    input [2:0] input_318;
    input [2:0] input_319;
    input [8:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      9'b000000000 : begin
        result = input_0;
      end
      9'b000000001 : begin
        result = input_1;
      end
      9'b000000010 : begin
        result = input_2;
      end
      9'b000000011 : begin
        result = input_3;
      end
      9'b000000100 : begin
        result = input_4;
      end
      9'b000000101 : begin
        result = input_5;
      end
      9'b000000110 : begin
        result = input_6;
      end
      9'b000000111 : begin
        result = input_7;
      end
      9'b000001000 : begin
        result = input_8;
      end
      9'b000001001 : begin
        result = input_9;
      end
      9'b000001010 : begin
        result = input_10;
      end
      9'b000001011 : begin
        result = input_11;
      end
      9'b000001100 : begin
        result = input_12;
      end
      9'b000001101 : begin
        result = input_13;
      end
      9'b000001110 : begin
        result = input_14;
      end
      9'b000001111 : begin
        result = input_15;
      end
      9'b000010000 : begin
        result = input_16;
      end
      9'b000010001 : begin
        result = input_17;
      end
      9'b000010010 : begin
        result = input_18;
      end
      9'b000010011 : begin
        result = input_19;
      end
      9'b000010100 : begin
        result = input_20;
      end
      9'b000010101 : begin
        result = input_21;
      end
      9'b000010110 : begin
        result = input_22;
      end
      9'b000010111 : begin
        result = input_23;
      end
      9'b000011000 : begin
        result = input_24;
      end
      9'b000011001 : begin
        result = input_25;
      end
      9'b000011010 : begin
        result = input_26;
      end
      9'b000011011 : begin
        result = input_27;
      end
      9'b000011100 : begin
        result = input_28;
      end
      9'b000011101 : begin
        result = input_29;
      end
      9'b000011110 : begin
        result = input_30;
      end
      9'b000011111 : begin
        result = input_31;
      end
      9'b000100000 : begin
        result = input_32;
      end
      9'b000100001 : begin
        result = input_33;
      end
      9'b000100010 : begin
        result = input_34;
      end
      9'b000100011 : begin
        result = input_35;
      end
      9'b000100100 : begin
        result = input_36;
      end
      9'b000100101 : begin
        result = input_37;
      end
      9'b000100110 : begin
        result = input_38;
      end
      9'b000100111 : begin
        result = input_39;
      end
      9'b000101000 : begin
        result = input_40;
      end
      9'b000101001 : begin
        result = input_41;
      end
      9'b000101010 : begin
        result = input_42;
      end
      9'b000101011 : begin
        result = input_43;
      end
      9'b000101100 : begin
        result = input_44;
      end
      9'b000101101 : begin
        result = input_45;
      end
      9'b000101110 : begin
        result = input_46;
      end
      9'b000101111 : begin
        result = input_47;
      end
      9'b000110000 : begin
        result = input_48;
      end
      9'b000110001 : begin
        result = input_49;
      end
      9'b000110010 : begin
        result = input_50;
      end
      9'b000110011 : begin
        result = input_51;
      end
      9'b000110100 : begin
        result = input_52;
      end
      9'b000110101 : begin
        result = input_53;
      end
      9'b000110110 : begin
        result = input_54;
      end
      9'b000110111 : begin
        result = input_55;
      end
      9'b000111000 : begin
        result = input_56;
      end
      9'b000111001 : begin
        result = input_57;
      end
      9'b000111010 : begin
        result = input_58;
      end
      9'b000111011 : begin
        result = input_59;
      end
      9'b000111100 : begin
        result = input_60;
      end
      9'b000111101 : begin
        result = input_61;
      end
      9'b000111110 : begin
        result = input_62;
      end
      9'b000111111 : begin
        result = input_63;
      end
      9'b001000000 : begin
        result = input_64;
      end
      9'b001000001 : begin
        result = input_65;
      end
      9'b001000010 : begin
        result = input_66;
      end
      9'b001000011 : begin
        result = input_67;
      end
      9'b001000100 : begin
        result = input_68;
      end
      9'b001000101 : begin
        result = input_69;
      end
      9'b001000110 : begin
        result = input_70;
      end
      9'b001000111 : begin
        result = input_71;
      end
      9'b001001000 : begin
        result = input_72;
      end
      9'b001001001 : begin
        result = input_73;
      end
      9'b001001010 : begin
        result = input_74;
      end
      9'b001001011 : begin
        result = input_75;
      end
      9'b001001100 : begin
        result = input_76;
      end
      9'b001001101 : begin
        result = input_77;
      end
      9'b001001110 : begin
        result = input_78;
      end
      9'b001001111 : begin
        result = input_79;
      end
      9'b001010000 : begin
        result = input_80;
      end
      9'b001010001 : begin
        result = input_81;
      end
      9'b001010010 : begin
        result = input_82;
      end
      9'b001010011 : begin
        result = input_83;
      end
      9'b001010100 : begin
        result = input_84;
      end
      9'b001010101 : begin
        result = input_85;
      end
      9'b001010110 : begin
        result = input_86;
      end
      9'b001010111 : begin
        result = input_87;
      end
      9'b001011000 : begin
        result = input_88;
      end
      9'b001011001 : begin
        result = input_89;
      end
      9'b001011010 : begin
        result = input_90;
      end
      9'b001011011 : begin
        result = input_91;
      end
      9'b001011100 : begin
        result = input_92;
      end
      9'b001011101 : begin
        result = input_93;
      end
      9'b001011110 : begin
        result = input_94;
      end
      9'b001011111 : begin
        result = input_95;
      end
      9'b001100000 : begin
        result = input_96;
      end
      9'b001100001 : begin
        result = input_97;
      end
      9'b001100010 : begin
        result = input_98;
      end
      9'b001100011 : begin
        result = input_99;
      end
      9'b001100100 : begin
        result = input_100;
      end
      9'b001100101 : begin
        result = input_101;
      end
      9'b001100110 : begin
        result = input_102;
      end
      9'b001100111 : begin
        result = input_103;
      end
      9'b001101000 : begin
        result = input_104;
      end
      9'b001101001 : begin
        result = input_105;
      end
      9'b001101010 : begin
        result = input_106;
      end
      9'b001101011 : begin
        result = input_107;
      end
      9'b001101100 : begin
        result = input_108;
      end
      9'b001101101 : begin
        result = input_109;
      end
      9'b001101110 : begin
        result = input_110;
      end
      9'b001101111 : begin
        result = input_111;
      end
      9'b001110000 : begin
        result = input_112;
      end
      9'b001110001 : begin
        result = input_113;
      end
      9'b001110010 : begin
        result = input_114;
      end
      9'b001110011 : begin
        result = input_115;
      end
      9'b001110100 : begin
        result = input_116;
      end
      9'b001110101 : begin
        result = input_117;
      end
      9'b001110110 : begin
        result = input_118;
      end
      9'b001110111 : begin
        result = input_119;
      end
      9'b001111000 : begin
        result = input_120;
      end
      9'b001111001 : begin
        result = input_121;
      end
      9'b001111010 : begin
        result = input_122;
      end
      9'b001111011 : begin
        result = input_123;
      end
      9'b001111100 : begin
        result = input_124;
      end
      9'b001111101 : begin
        result = input_125;
      end
      9'b001111110 : begin
        result = input_126;
      end
      9'b001111111 : begin
        result = input_127;
      end
      9'b010000000 : begin
        result = input_128;
      end
      9'b010000001 : begin
        result = input_129;
      end
      9'b010000010 : begin
        result = input_130;
      end
      9'b010000011 : begin
        result = input_131;
      end
      9'b010000100 : begin
        result = input_132;
      end
      9'b010000101 : begin
        result = input_133;
      end
      9'b010000110 : begin
        result = input_134;
      end
      9'b010000111 : begin
        result = input_135;
      end
      9'b010001000 : begin
        result = input_136;
      end
      9'b010001001 : begin
        result = input_137;
      end
      9'b010001010 : begin
        result = input_138;
      end
      9'b010001011 : begin
        result = input_139;
      end
      9'b010001100 : begin
        result = input_140;
      end
      9'b010001101 : begin
        result = input_141;
      end
      9'b010001110 : begin
        result = input_142;
      end
      9'b010001111 : begin
        result = input_143;
      end
      9'b010010000 : begin
        result = input_144;
      end
      9'b010010001 : begin
        result = input_145;
      end
      9'b010010010 : begin
        result = input_146;
      end
      9'b010010011 : begin
        result = input_147;
      end
      9'b010010100 : begin
        result = input_148;
      end
      9'b010010101 : begin
        result = input_149;
      end
      9'b010010110 : begin
        result = input_150;
      end
      9'b010010111 : begin
        result = input_151;
      end
      9'b010011000 : begin
        result = input_152;
      end
      9'b010011001 : begin
        result = input_153;
      end
      9'b010011010 : begin
        result = input_154;
      end
      9'b010011011 : begin
        result = input_155;
      end
      9'b010011100 : begin
        result = input_156;
      end
      9'b010011101 : begin
        result = input_157;
      end
      9'b010011110 : begin
        result = input_158;
      end
      9'b010011111 : begin
        result = input_159;
      end
      9'b010100000 : begin
        result = input_160;
      end
      9'b010100001 : begin
        result = input_161;
      end
      9'b010100010 : begin
        result = input_162;
      end
      9'b010100011 : begin
        result = input_163;
      end
      9'b010100100 : begin
        result = input_164;
      end
      9'b010100101 : begin
        result = input_165;
      end
      9'b010100110 : begin
        result = input_166;
      end
      9'b010100111 : begin
        result = input_167;
      end
      9'b010101000 : begin
        result = input_168;
      end
      9'b010101001 : begin
        result = input_169;
      end
      9'b010101010 : begin
        result = input_170;
      end
      9'b010101011 : begin
        result = input_171;
      end
      9'b010101100 : begin
        result = input_172;
      end
      9'b010101101 : begin
        result = input_173;
      end
      9'b010101110 : begin
        result = input_174;
      end
      9'b010101111 : begin
        result = input_175;
      end
      9'b010110000 : begin
        result = input_176;
      end
      9'b010110001 : begin
        result = input_177;
      end
      9'b010110010 : begin
        result = input_178;
      end
      9'b010110011 : begin
        result = input_179;
      end
      9'b010110100 : begin
        result = input_180;
      end
      9'b010110101 : begin
        result = input_181;
      end
      9'b010110110 : begin
        result = input_182;
      end
      9'b010110111 : begin
        result = input_183;
      end
      9'b010111000 : begin
        result = input_184;
      end
      9'b010111001 : begin
        result = input_185;
      end
      9'b010111010 : begin
        result = input_186;
      end
      9'b010111011 : begin
        result = input_187;
      end
      9'b010111100 : begin
        result = input_188;
      end
      9'b010111101 : begin
        result = input_189;
      end
      9'b010111110 : begin
        result = input_190;
      end
      9'b010111111 : begin
        result = input_191;
      end
      9'b011000000 : begin
        result = input_192;
      end
      9'b011000001 : begin
        result = input_193;
      end
      9'b011000010 : begin
        result = input_194;
      end
      9'b011000011 : begin
        result = input_195;
      end
      9'b011000100 : begin
        result = input_196;
      end
      9'b011000101 : begin
        result = input_197;
      end
      9'b011000110 : begin
        result = input_198;
      end
      9'b011000111 : begin
        result = input_199;
      end
      9'b011001000 : begin
        result = input_200;
      end
      9'b011001001 : begin
        result = input_201;
      end
      9'b011001010 : begin
        result = input_202;
      end
      9'b011001011 : begin
        result = input_203;
      end
      9'b011001100 : begin
        result = input_204;
      end
      9'b011001101 : begin
        result = input_205;
      end
      9'b011001110 : begin
        result = input_206;
      end
      9'b011001111 : begin
        result = input_207;
      end
      9'b011010000 : begin
        result = input_208;
      end
      9'b011010001 : begin
        result = input_209;
      end
      9'b011010010 : begin
        result = input_210;
      end
      9'b011010011 : begin
        result = input_211;
      end
      9'b011010100 : begin
        result = input_212;
      end
      9'b011010101 : begin
        result = input_213;
      end
      9'b011010110 : begin
        result = input_214;
      end
      9'b011010111 : begin
        result = input_215;
      end
      9'b011011000 : begin
        result = input_216;
      end
      9'b011011001 : begin
        result = input_217;
      end
      9'b011011010 : begin
        result = input_218;
      end
      9'b011011011 : begin
        result = input_219;
      end
      9'b011011100 : begin
        result = input_220;
      end
      9'b011011101 : begin
        result = input_221;
      end
      9'b011011110 : begin
        result = input_222;
      end
      9'b011011111 : begin
        result = input_223;
      end
      9'b011100000 : begin
        result = input_224;
      end
      9'b011100001 : begin
        result = input_225;
      end
      9'b011100010 : begin
        result = input_226;
      end
      9'b011100011 : begin
        result = input_227;
      end
      9'b011100100 : begin
        result = input_228;
      end
      9'b011100101 : begin
        result = input_229;
      end
      9'b011100110 : begin
        result = input_230;
      end
      9'b011100111 : begin
        result = input_231;
      end
      9'b011101000 : begin
        result = input_232;
      end
      9'b011101001 : begin
        result = input_233;
      end
      9'b011101010 : begin
        result = input_234;
      end
      9'b011101011 : begin
        result = input_235;
      end
      9'b011101100 : begin
        result = input_236;
      end
      9'b011101101 : begin
        result = input_237;
      end
      9'b011101110 : begin
        result = input_238;
      end
      9'b011101111 : begin
        result = input_239;
      end
      9'b011110000 : begin
        result = input_240;
      end
      9'b011110001 : begin
        result = input_241;
      end
      9'b011110010 : begin
        result = input_242;
      end
      9'b011110011 : begin
        result = input_243;
      end
      9'b011110100 : begin
        result = input_244;
      end
      9'b011110101 : begin
        result = input_245;
      end
      9'b011110110 : begin
        result = input_246;
      end
      9'b011110111 : begin
        result = input_247;
      end
      9'b011111000 : begin
        result = input_248;
      end
      9'b011111001 : begin
        result = input_249;
      end
      9'b011111010 : begin
        result = input_250;
      end
      9'b011111011 : begin
        result = input_251;
      end
      9'b011111100 : begin
        result = input_252;
      end
      9'b011111101 : begin
        result = input_253;
      end
      9'b011111110 : begin
        result = input_254;
      end
      9'b011111111 : begin
        result = input_255;
      end
      9'b100000000 : begin
        result = input_256;
      end
      9'b100000001 : begin
        result = input_257;
      end
      9'b100000010 : begin
        result = input_258;
      end
      9'b100000011 : begin
        result = input_259;
      end
      9'b100000100 : begin
        result = input_260;
      end
      9'b100000101 : begin
        result = input_261;
      end
      9'b100000110 : begin
        result = input_262;
      end
      9'b100000111 : begin
        result = input_263;
      end
      9'b100001000 : begin
        result = input_264;
      end
      9'b100001001 : begin
        result = input_265;
      end
      9'b100001010 : begin
        result = input_266;
      end
      9'b100001011 : begin
        result = input_267;
      end
      9'b100001100 : begin
        result = input_268;
      end
      9'b100001101 : begin
        result = input_269;
      end
      9'b100001110 : begin
        result = input_270;
      end
      9'b100001111 : begin
        result = input_271;
      end
      9'b100010000 : begin
        result = input_272;
      end
      9'b100010001 : begin
        result = input_273;
      end
      9'b100010010 : begin
        result = input_274;
      end
      9'b100010011 : begin
        result = input_275;
      end
      9'b100010100 : begin
        result = input_276;
      end
      9'b100010101 : begin
        result = input_277;
      end
      9'b100010110 : begin
        result = input_278;
      end
      9'b100010111 : begin
        result = input_279;
      end
      9'b100011000 : begin
        result = input_280;
      end
      9'b100011001 : begin
        result = input_281;
      end
      9'b100011010 : begin
        result = input_282;
      end
      9'b100011011 : begin
        result = input_283;
      end
      9'b100011100 : begin
        result = input_284;
      end
      9'b100011101 : begin
        result = input_285;
      end
      9'b100011110 : begin
        result = input_286;
      end
      9'b100011111 : begin
        result = input_287;
      end
      9'b100100000 : begin
        result = input_288;
      end
      9'b100100001 : begin
        result = input_289;
      end
      9'b100100010 : begin
        result = input_290;
      end
      9'b100100011 : begin
        result = input_291;
      end
      9'b100100100 : begin
        result = input_292;
      end
      9'b100100101 : begin
        result = input_293;
      end
      9'b100100110 : begin
        result = input_294;
      end
      9'b100100111 : begin
        result = input_295;
      end
      9'b100101000 : begin
        result = input_296;
      end
      9'b100101001 : begin
        result = input_297;
      end
      9'b100101010 : begin
        result = input_298;
      end
      9'b100101011 : begin
        result = input_299;
      end
      9'b100101100 : begin
        result = input_300;
      end
      9'b100101101 : begin
        result = input_301;
      end
      9'b100101110 : begin
        result = input_302;
      end
      9'b100101111 : begin
        result = input_303;
      end
      9'b100110000 : begin
        result = input_304;
      end
      9'b100110001 : begin
        result = input_305;
      end
      9'b100110010 : begin
        result = input_306;
      end
      9'b100110011 : begin
        result = input_307;
      end
      9'b100110100 : begin
        result = input_308;
      end
      9'b100110101 : begin
        result = input_309;
      end
      9'b100110110 : begin
        result = input_310;
      end
      9'b100110111 : begin
        result = input_311;
      end
      9'b100111000 : begin
        result = input_312;
      end
      9'b100111001 : begin
        result = input_313;
      end
      9'b100111010 : begin
        result = input_314;
      end
      9'b100111011 : begin
        result = input_315;
      end
      9'b100111100 : begin
        result = input_316;
      end
      9'b100111101 : begin
        result = input_317;
      end
      9'b100111110 : begin
        result = input_318;
      end
      default : begin
        result = input_319;
      end
    endcase
    MUX_v_3_320_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i3_1o8_b7f1baaf117249900fa3606aa9bde444b0_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Fri Nov  1 23:14:08 2019
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i3_1o8_b7f1baaf117249900fa3606aa9bde444b0
// ------------------------------------------------------------------


module ROM_1i3_1o8_b7f1baaf117249900fa3606aa9bde444b0 (
  I_1, O_1
);
  input [2:0] I_1;
  output [7:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_8_8_2(8'b00011100, 8'b01001011, 8'b01101100, 8'b10000100, 8'b10010111,
      8'b10100110, 8'b10110011, 8'b10111100, I_1);

  function automatic [7:0] MUX_v_8_8_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [2:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_8_8_2 = result;
  end
  endfunction

endmodule




//------> /opt/cad/catapult/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ../td_ccore_solutions/leading_sign_71_0_e5d4bd9dc928fda5adf5bf26ec9a2550b9a2_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Fri Nov  1 23:14:19 2019
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_71_0
// ------------------------------------------------------------------


module leading_sign_71_0 (
  mantissa, rtn
);
  input [70:0] mantissa;
  output [6:0] rtn;


  // Interconnect Declarations
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_6_2_sdt_2;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_18_3_sdt_3;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_26_2_sdt_2;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_42_4_sdt_4;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_50_2_sdt_2;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_62_3_sdt_3;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_70_2_sdt_2;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_90_5_sdt_5;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_98_2_sdt_2;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_110_3_sdt_3;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_118_2_sdt_2;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_134_4_sdt_4;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_142_2_sdt_2;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_154_3_sdt_3;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_162_2_sdt_2;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_186_6_sdt_6;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_194_2_sdt_2;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_6_2_sdt_1;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_14_2_sdt_1;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_26_2_sdt_1;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_34_2_sdt_1;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_50_2_sdt_1;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_58_2_sdt_1;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_70_2_sdt_1;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_78_2_sdt_1;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_98_2_sdt_1;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_106_2_sdt_1;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_118_2_sdt_1;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_126_2_sdt_1;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_142_2_sdt_1;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_150_2_sdt_1;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_162_2_sdt_1;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_170_2_sdt_1;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_194_2_sdt_1;
  wire ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_200_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;
  wire c_h_1_17;
  wire c_h_1_20;
  wire c_h_1_21;
  wire c_h_1_24;
  wire c_h_1_27;
  wire c_h_1_28;
  wire c_h_1_29;
  wire c_h_1_30;
  wire c_h_1_33;
  wire c_h_1_34;

  wire[0:0] ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_nl;
  wire[0:0] ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_1_nl;
  wire[0:0] ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_2_nl;
  wire[2:0] ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_or_1_nl;
  wire[0:0] ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_293_nl;
  wire[0:0] ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_295_nl;
  wire[0:0] ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_296_nl;
  wire[0:0] ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_281_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_6_2_sdt_2
      = ~((mantissa[68:67]!=2'b00));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_6_2_sdt_1
      = ~((mantissa[70:69]!=2'b00));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_14_2_sdt_1
      = ~((mantissa[66:65]!=2'b00));
  assign c_h_1_2 = ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_6_2_sdt_1
      & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_6_2_sdt_2;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_18_3_sdt_3
      = (mantissa[64:63]==2'b00) & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_14_2_sdt_1;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_26_2_sdt_2
      = ~((mantissa[60:59]!=2'b00));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_26_2_sdt_1
      = ~((mantissa[62:61]!=2'b00));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_34_2_sdt_1
      = ~((mantissa[58:57]!=2'b00));
  assign c_h_1_5 = ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_26_2_sdt_1
      & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_18_3_sdt_3;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_42_4_sdt_4
      = (mantissa[56:55]==2'b00) & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_34_2_sdt_1
      & c_h_1_5;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_50_2_sdt_2
      = ~((mantissa[52:51]!=2'b00));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_50_2_sdt_1
      = ~((mantissa[54:53]!=2'b00));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_58_2_sdt_1
      = ~((mantissa[50:49]!=2'b00));
  assign c_h_1_9 = ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_50_2_sdt_1
      & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_50_2_sdt_2;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_62_3_sdt_3
      = (mantissa[48:47]==2'b00) & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_58_2_sdt_1;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_70_2_sdt_2
      = ~((mantissa[44:43]!=2'b00));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_70_2_sdt_1
      = ~((mantissa[46:45]!=2'b00));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_78_2_sdt_1
      = ~((mantissa[42:41]!=2'b00));
  assign c_h_1_12 = ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_70_2_sdt_1
      & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_42_4_sdt_4;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_90_5_sdt_5
      = (mantissa[40:39]==2'b00) & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_78_2_sdt_1
      & c_h_1_12 & c_h_1_13;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_98_2_sdt_2
      = ~((mantissa[36:35]!=2'b00));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_98_2_sdt_1
      = ~((mantissa[38:37]!=2'b00));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_106_2_sdt_1
      = ~((mantissa[34:33]!=2'b00));
  assign c_h_1_17 = ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_98_2_sdt_1
      & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_98_2_sdt_2;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_110_3_sdt_3
      = (mantissa[32:31]==2'b00) & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_106_2_sdt_1;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_118_2_sdt_2
      = ~((mantissa[28:27]!=2'b00));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_118_2_sdt_1
      = ~((mantissa[30:29]!=2'b00));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_126_2_sdt_1
      = ~((mantissa[26:25]!=2'b00));
  assign c_h_1_20 = ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_118_2_sdt_1
      & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_118_2_sdt_2;
  assign c_h_1_21 = c_h_1_17 & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_110_3_sdt_3;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_134_4_sdt_4
      = (mantissa[24:23]==2'b00) & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_126_2_sdt_1
      & c_h_1_20;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_142_2_sdt_2
      = ~((mantissa[20:19]!=2'b00));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_142_2_sdt_1
      = ~((mantissa[22:21]!=2'b00));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_150_2_sdt_1
      = ~((mantissa[18:17]!=2'b00));
  assign c_h_1_24 = ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_142_2_sdt_1
      & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_142_2_sdt_2;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_154_3_sdt_3
      = (mantissa[16:15]==2'b00) & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_150_2_sdt_1;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_162_2_sdt_2
      = ~((mantissa[12:11]!=2'b00));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_162_2_sdt_1
      = ~((mantissa[14:13]!=2'b00));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_170_2_sdt_1
      = ~((mantissa[10:9]!=2'b00));
  assign c_h_1_27 = ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_162_2_sdt_1
      & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_162_2_sdt_2;
  assign c_h_1_28 = c_h_1_24 & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_154_3_sdt_3;
  assign c_h_1_29 = c_h_1_21 & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_134_4_sdt_4;
  assign c_h_1_30 = c_h_1_14 & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_90_5_sdt_5;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_186_6_sdt_6
      = (mantissa[8:7]==2'b00) & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_170_2_sdt_1
      & c_h_1_27 & c_h_1_28 & c_h_1_29;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_194_2_sdt_2
      = ~((mantissa[4:3]!=2'b00));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_194_2_sdt_1
      = ~((mantissa[6:5]!=2'b00));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_200_2_sdt_1
      = ~((mantissa[2:1]!=2'b00));
  assign c_h_1_33 = ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_194_2_sdt_1
      & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_194_2_sdt_2;
  assign c_h_1_34 = c_h_1_30 & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_186_6_sdt_6;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_nl
      = c_h_1_30 & (~ ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_186_6_sdt_6);
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_1_nl
      = c_h_1_14 & (c_h_1_29 | (~ ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_90_5_sdt_5))
      & (~ c_h_1_34);
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_2_nl
      = c_h_1_6 & (c_h_1_13 | (~ ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_42_4_sdt_4))
      & (~((~(c_h_1_21 & (c_h_1_28 | (~ ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_134_4_sdt_4))))
      & c_h_1_30)) & (~ c_h_1_34);
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_293_nl
      = c_h_1_2 & (c_h_1_5 | (~ ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_18_3_sdt_3))
      & (~((~(c_h_1_9 & (c_h_1_12 | (~ ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_62_3_sdt_3))))
      & c_h_1_14)) & (~((~(c_h_1_17 & (c_h_1_20 | (~ ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_110_3_sdt_3))
      & (~((~(c_h_1_24 & (c_h_1_27 | (~ ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_154_3_sdt_3))))
      & c_h_1_29)))) & c_h_1_30)) & (c_h_1_33 | (~ c_h_1_34));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_295_nl
      = ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_6_2_sdt_1
      & (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_14_2_sdt_1
      | (~ ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_26_2_sdt_1
      & (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_34_2_sdt_1
      | (~ ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_26_2_sdt_2))))
      & c_h_1_6)) & (~((~(ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_50_2_sdt_1
      & (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_58_2_sdt_1
      | (~ ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_50_2_sdt_2))
      & (~((~(ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_70_2_sdt_1
      & (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_78_2_sdt_1
      | (~ ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14)) & (~((~(ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_98_2_sdt_1
      & (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_106_2_sdt_1
      | (~ ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_98_2_sdt_2))
      & (~((~(ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_118_2_sdt_1
      & (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_126_2_sdt_1
      | (~ ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_118_2_sdt_2))))
      & c_h_1_21)) & (~((~(ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_142_2_sdt_1
      & (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_150_2_sdt_1
      | (~ ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_142_2_sdt_2))
      & (~((~(ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_162_2_sdt_1
      & (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_170_2_sdt_1
      | (~ ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_162_2_sdt_2))))
      & c_h_1_28)))) & c_h_1_29)))) & c_h_1_30)) & (~((~(ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_194_2_sdt_1
      & (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_200_2_sdt_1
      | (~ ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_194_2_sdt_2))))
      & c_h_1_34));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_296_nl
      = (~((mantissa[70]) | (~((mantissa[69:68]!=2'b01))))) & (~(((mantissa[66])
      | (~((mantissa[65:64]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[62]) | (~((mantissa[61:60]!=2'b01)))))
      & (~(((mantissa[58]) | (~((mantissa[57:56]!=2'b01)))) & c_h_1_5)))) & c_h_1_6))
      & (~((~((~((mantissa[54]) | (~((mantissa[53:52]!=2'b01))))) & (~(((mantissa[50])
      | (~((mantissa[49:48]!=2'b01)))) & c_h_1_9)) & (~((~((~((mantissa[46]) | (~((mantissa[45:44]!=2'b01)))))
      & (~(((mantissa[42]) | (~((mantissa[41:40]!=2'b01)))) & c_h_1_12)))) & c_h_1_13))))
      & c_h_1_14)) & (~((~((~((mantissa[38]) | (~((mantissa[37:36]!=2'b01))))) &
      (~(((mantissa[34]) | (~((mantissa[33:32]!=2'b01)))) & c_h_1_17)) & (~((~((~((mantissa[30])
      | (~((mantissa[29:28]!=2'b01))))) & (~(((mantissa[26]) | (~((mantissa[25:24]!=2'b01))))
      & c_h_1_20)))) & c_h_1_21)) & (~((~((~((mantissa[22]) | (~((mantissa[21:20]!=2'b01)))))
      & (~(((mantissa[18]) | (~((mantissa[17:16]!=2'b01)))) & c_h_1_24)) & (~((~((~((mantissa[14])
      | (~((mantissa[13:12]!=2'b01))))) & (~(((mantissa[10]) | (~((mantissa[9:8]!=2'b01))))
      & c_h_1_27)))) & c_h_1_28)))) & c_h_1_29)))) & c_h_1_30)) & (~((~((~((mantissa[6])
      | (~((mantissa[5:4]!=2'b01))))) & (~((~((mantissa[2:1]==2'b01))) & c_h_1_33))))
      & c_h_1_34));
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_281_nl
      = (~ (mantissa[0])) & ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_wrs_c_200_2_sdt_1
      & c_h_1_33 & c_h_1_34;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_or_1_nl
      = MUX_v_3_2_2(({(ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_293_nl)
      , (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_295_nl)
      , (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_296_nl)}),
      3'b111, (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_281_nl));
  assign rtn = {c_h_1_34 , (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_nl)
      , (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_1_nl)
      , (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_and_2_nl)
      , (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_leading_1_leading_sign_71_0_rtn_or_1_nl)};

  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction

endmodule




//------> /opt/cad/catapult/pkgs/siflibs/mgc_shift_bl_beh_v5.v 
module mgc_shift_bl_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate if ( signd_a )
   begin: SGNED
     assign z = fshl_s(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
     assign z = fshl_s(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift left - signed shift argument
   function [width_z-1:0] fshl_s;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      reg [width_a:0] sbit_arg1;
      begin
        // Ignoring the possibility that arg2[width_s-1] could be X
        // because of customer complaints regarding X'es in simulation results
        if ( arg2[width_s-1] == 1'b0 )
        begin
          sbit_arg1[width_a:0] = {(width_a+1){1'b0}};
          fshl_s = fshl_u(arg1, arg2, sbit);
        end
        else
        begin
          sbit_arg1[width_a] = sbit;
          sbit_arg1[width_a-1:0] = arg1;
          fshl_s = fshr_u(sbit_arg1[width_a:1], ~arg2, sbit);
        end
      end
   endfunction

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Sat Nov  2 11:12:10 2019
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_ccs_sample_mem_ccs_ram_sync_dualport_rwport_9_18_10_640_640_18_5_gen
// ------------------------------------------------------------------


module mnist_mlp_ccs_sample_mem_ccs_ram_sync_dualport_rwport_9_18_10_640_640_18_5_gen
    (
  qb, web, enb, db, adrb, qa, wea, ena, da, adra, adra_d, da_d, ena_d, wea_d, qa_d,
      port_0_rw_ram_ir_internal_RMASK_B_d, port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [17:0] qb;
  output web;
  output enb;
  output [17:0] db;
  output [9:0] adrb;
  input [17:0] qa;
  output wea;
  output ena;
  output [17:0] da;
  output [9:0] adra;
  input [19:0] adra_d;
  input [35:0] da_d;
  input [1:0] ena_d;
  input [1:0] wea_d;
  output [35:0] qa_d;
  input [1:0] port_0_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] port_0_rw_ram_ir_internal_WMASK_B_d;


  wire w6_or_nl;
  wire w6_or_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign qa_d[35:18] = qb;
  assign web = (port_0_rw_ram_ir_internal_WMASK_B_d[1]);
  assign w6_or_nl = (port_0_rw_ram_ir_internal_RMASK_B_d[1]) | (port_0_rw_ram_ir_internal_WMASK_B_d[1]);
  assign enb = (w6_or_nl);
  assign db = (da_d[35:18]);
  assign adrb = (adra_d[19:10]);
  assign qa_d[17:0] = qa;
  assign wea = (port_0_rw_ram_ir_internal_WMASK_B_d[0]);
  assign w6_or_1_nl = (port_0_rw_ram_ir_internal_RMASK_B_d[0]) | (port_0_rw_ram_ir_internal_WMASK_B_d[0]);
  assign ena = (w6_or_1_nl);
  assign da = (da_d[17:0]);
  assign adra = (adra_d[9:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_ccs_sample_mem_ccs_ram_sync_dualport_rwport_7_18_12_4096_4096_18_5_gen
// ------------------------------------------------------------------


module mnist_mlp_ccs_sample_mem_ccs_ram_sync_dualport_rwport_7_18_12_4096_4096_18_5_gen
    (
  qb, web, enb, db, adrb, qa, wea, ena, da, adra, adra_d, da_d, ena_d, wea_d, qa_d,
      port_0_rw_ram_ir_internal_RMASK_B_d, port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [17:0] qb;
  output web;
  output enb;
  output [17:0] db;
  output [11:0] adrb;
  input [17:0] qa;
  output wea;
  output ena;
  output [17:0] da;
  output [11:0] adra;
  input [23:0] adra_d;
  input [35:0] da_d;
  input [1:0] ena_d;
  input [1:0] wea_d;
  output [35:0] qa_d;
  input [1:0] port_0_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] port_0_rw_ram_ir_internal_WMASK_B_d;


  wire w4_or_nl;
  wire w4_or_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign qa_d[35:18] = qb;
  assign web = (port_0_rw_ram_ir_internal_WMASK_B_d[1]);
  assign w4_or_nl = (port_0_rw_ram_ir_internal_RMASK_B_d[1]) | (port_0_rw_ram_ir_internal_WMASK_B_d[1]);
  assign enb = (w4_or_nl);
  assign db = (da_d[35:18]);
  assign adrb = (adra_d[23:12]);
  assign qa_d[17:0] = qa;
  assign wea = (port_0_rw_ram_ir_internal_WMASK_B_d[0]);
  assign w4_or_1_nl = (port_0_rw_ram_ir_internal_RMASK_B_d[0]) | (port_0_rw_ram_ir_internal_WMASK_B_d[0]);
  assign ena = (w4_or_1_nl);
  assign da = (da_d[17:0]);
  assign adra = (adra_d[11:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_ccs_sample_mem_ccs_ram_sync_dualport_rwport_5_18_16_50176_50176_18_5_gen
// ------------------------------------------------------------------


module mnist_mlp_ccs_sample_mem_ccs_ram_sync_dualport_rwport_5_18_16_50176_50176_18_5_gen
    (
  qb, web, enb, db, adrb, qa, wea, ena, da, adra, adra_d, da_d, ena_d, wea_d, qa_d,
      port_0_rw_ram_ir_internal_RMASK_B_d, port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [17:0] qb;
  output web;
  output enb;
  output [17:0] db;
  output [15:0] adrb;
  input [17:0] qa;
  output wea;
  output ena;
  output [17:0] da;
  output [15:0] adra;
  input [31:0] adra_d;
  input [35:0] da_d;
  input [1:0] ena_d;
  input [1:0] wea_d;
  output [35:0] qa_d;
  input [1:0] port_0_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] port_0_rw_ram_ir_internal_WMASK_B_d;


  wire w2_or_nl;
  wire w2_or_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign qa_d[35:18] = qb;
  assign web = (port_0_rw_ram_ir_internal_WMASK_B_d[1]);
  assign w2_or_nl = (port_0_rw_ram_ir_internal_RMASK_B_d[1]) | (port_0_rw_ram_ir_internal_WMASK_B_d[1]);
  assign enb = (w2_or_nl);
  assign db = (da_d[35:18]);
  assign adrb = (adra_d[31:16]);
  assign qa_d[17:0] = qa;
  assign wea = (port_0_rw_ram_ir_internal_WMASK_B_d[0]);
  assign w2_or_1_nl = (port_0_rw_ram_ir_internal_RMASK_B_d[0]) | (port_0_rw_ram_ir_internal_WMASK_B_d[0]);
  assign ena = (w2_or_1_nl);
  assign da = (da_d[17:0]);
  assign adra = (adra_d[15:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module mnist_mlp_core_core_fsm (
  clk, rst, core_wen, fsm_output, InitAccumLoop_C_0_tr0, IndexLoop_C_0_tr0, InitAccumLoop_1_C_0_tr0,
      ReuseLoop_1_C_0_tr0, InitAccumLoop_2_C_0_tr0, ReuseLoop_2_C_0_tr0, nnet_softmax_layer6_t_result_t_softmax_config7_for_1_C_0_tr0
);
  input clk;
  input rst;
  input core_wen;
  output [7:0] fsm_output;
  reg [7:0] fsm_output;
  input InitAccumLoop_C_0_tr0;
  input IndexLoop_C_0_tr0;
  input InitAccumLoop_1_C_0_tr0;
  input ReuseLoop_1_C_0_tr0;
  input InitAccumLoop_2_C_0_tr0;
  input ReuseLoop_2_C_0_tr0;
  input nnet_softmax_layer6_t_result_t_softmax_config7_for_1_C_0_tr0;


  // FSM State Type Declaration for mnist_mlp_core_core_fsm_1
  parameter
    core_rlp_C_0 = 8'd0,
    main_C_0 = 8'd1,
    InitAccumLoop_C_0 = 8'd2,
    IndexLoop_C_0 = 8'd3,
    main_C_1 = 8'd4,
    main_C_2 = 8'd5,
    main_C_3 = 8'd6,
    main_C_4 = 8'd7,
    main_C_5 = 8'd8,
    main_C_6 = 8'd9,
    main_C_7 = 8'd10,
    main_C_8 = 8'd11,
    main_C_9 = 8'd12,
    main_C_10 = 8'd13,
    main_C_11 = 8'd14,
    main_C_12 = 8'd15,
    main_C_13 = 8'd16,
    main_C_14 = 8'd17,
    main_C_15 = 8'd18,
    main_C_16 = 8'd19,
    main_C_17 = 8'd20,
    main_C_18 = 8'd21,
    main_C_19 = 8'd22,
    main_C_20 = 8'd23,
    main_C_21 = 8'd24,
    main_C_22 = 8'd25,
    main_C_23 = 8'd26,
    main_C_24 = 8'd27,
    main_C_25 = 8'd28,
    main_C_26 = 8'd29,
    main_C_27 = 8'd30,
    main_C_28 = 8'd31,
    main_C_29 = 8'd32,
    main_C_30 = 8'd33,
    main_C_31 = 8'd34,
    main_C_32 = 8'd35,
    main_C_33 = 8'd36,
    main_C_34 = 8'd37,
    main_C_35 = 8'd38,
    main_C_36 = 8'd39,
    main_C_37 = 8'd40,
    main_C_38 = 8'd41,
    main_C_39 = 8'd42,
    main_C_40 = 8'd43,
    main_C_41 = 8'd44,
    main_C_42 = 8'd45,
    main_C_43 = 8'd46,
    main_C_44 = 8'd47,
    main_C_45 = 8'd48,
    main_C_46 = 8'd49,
    main_C_47 = 8'd50,
    main_C_48 = 8'd51,
    main_C_49 = 8'd52,
    main_C_50 = 8'd53,
    main_C_51 = 8'd54,
    main_C_52 = 8'd55,
    main_C_53 = 8'd56,
    main_C_54 = 8'd57,
    main_C_55 = 8'd58,
    main_C_56 = 8'd59,
    main_C_57 = 8'd60,
    main_C_58 = 8'd61,
    main_C_59 = 8'd62,
    main_C_60 = 8'd63,
    main_C_61 = 8'd64,
    main_C_62 = 8'd65,
    main_C_63 = 8'd66,
    main_C_64 = 8'd67,
    InitAccumLoop_1_C_0 = 8'd68,
    ReuseLoop_1_C_0 = 8'd69,
    main_C_65 = 8'd70,
    main_C_66 = 8'd71,
    main_C_67 = 8'd72,
    main_C_68 = 8'd73,
    main_C_69 = 8'd74,
    main_C_70 = 8'd75,
    main_C_71 = 8'd76,
    main_C_72 = 8'd77,
    main_C_73 = 8'd78,
    main_C_74 = 8'd79,
    main_C_75 = 8'd80,
    main_C_76 = 8'd81,
    main_C_77 = 8'd82,
    main_C_78 = 8'd83,
    main_C_79 = 8'd84,
    main_C_80 = 8'd85,
    main_C_81 = 8'd86,
    main_C_82 = 8'd87,
    main_C_83 = 8'd88,
    main_C_84 = 8'd89,
    main_C_85 = 8'd90,
    main_C_86 = 8'd91,
    main_C_87 = 8'd92,
    main_C_88 = 8'd93,
    main_C_89 = 8'd94,
    main_C_90 = 8'd95,
    main_C_91 = 8'd96,
    main_C_92 = 8'd97,
    main_C_93 = 8'd98,
    main_C_94 = 8'd99,
    main_C_95 = 8'd100,
    main_C_96 = 8'd101,
    main_C_97 = 8'd102,
    main_C_98 = 8'd103,
    main_C_99 = 8'd104,
    main_C_100 = 8'd105,
    main_C_101 = 8'd106,
    main_C_102 = 8'd107,
    main_C_103 = 8'd108,
    main_C_104 = 8'd109,
    main_C_105 = 8'd110,
    main_C_106 = 8'd111,
    main_C_107 = 8'd112,
    main_C_108 = 8'd113,
    main_C_109 = 8'd114,
    main_C_110 = 8'd115,
    main_C_111 = 8'd116,
    main_C_112 = 8'd117,
    main_C_113 = 8'd118,
    main_C_114 = 8'd119,
    main_C_115 = 8'd120,
    main_C_116 = 8'd121,
    main_C_117 = 8'd122,
    main_C_118 = 8'd123,
    main_C_119 = 8'd124,
    main_C_120 = 8'd125,
    main_C_121 = 8'd126,
    main_C_122 = 8'd127,
    main_C_123 = 8'd128,
    main_C_124 = 8'd129,
    main_C_125 = 8'd130,
    main_C_126 = 8'd131,
    main_C_127 = 8'd132,
    main_C_128 = 8'd133,
    InitAccumLoop_2_C_0 = 8'd134,
    ReuseLoop_2_C_0 = 8'd135,
    main_C_129 = 8'd136,
    main_C_130 = 8'd137,
    main_C_131 = 8'd138,
    main_C_132 = 8'd139,
    main_C_133 = 8'd140,
    main_C_134 = 8'd141,
    main_C_135 = 8'd142,
    main_C_136 = 8'd143,
    main_C_137 = 8'd144,
    main_C_138 = 8'd145,
    main_C_139 = 8'd146,
    main_C_140 = 8'd147,
    main_C_141 = 8'd148,
    main_C_142 = 8'd149,
    main_C_143 = 8'd150,
    main_C_144 = 8'd151,
    main_C_145 = 8'd152,
    main_C_146 = 8'd153,
    main_C_147 = 8'd154,
    main_C_148 = 8'd155,
    main_C_149 = 8'd156,
    main_C_150 = 8'd157,
    nnet_softmax_layer6_t_result_t_softmax_config7_for_1_C_0 = 8'd158;

  reg [7:0] state_var;
  reg [7:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : mnist_mlp_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 8'b00000001;
        state_var_NS = InitAccumLoop_C_0;
      end
      InitAccumLoop_C_0 : begin
        fsm_output = 8'b00000010;
        if ( InitAccumLoop_C_0_tr0 ) begin
          state_var_NS = IndexLoop_C_0;
        end
        else begin
          state_var_NS = InitAccumLoop_C_0;
        end
      end
      IndexLoop_C_0 : begin
        fsm_output = 8'b00000011;
        if ( IndexLoop_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = IndexLoop_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 8'b00000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 8'b00000101;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 8'b00000110;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 8'b00000111;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 8'b00001000;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 8'b00001001;
        state_var_NS = main_C_7;
      end
      main_C_7 : begin
        fsm_output = 8'b00001010;
        state_var_NS = main_C_8;
      end
      main_C_8 : begin
        fsm_output = 8'b00001011;
        state_var_NS = main_C_9;
      end
      main_C_9 : begin
        fsm_output = 8'b00001100;
        state_var_NS = main_C_10;
      end
      main_C_10 : begin
        fsm_output = 8'b00001101;
        state_var_NS = main_C_11;
      end
      main_C_11 : begin
        fsm_output = 8'b00001110;
        state_var_NS = main_C_12;
      end
      main_C_12 : begin
        fsm_output = 8'b00001111;
        state_var_NS = main_C_13;
      end
      main_C_13 : begin
        fsm_output = 8'b00010000;
        state_var_NS = main_C_14;
      end
      main_C_14 : begin
        fsm_output = 8'b00010001;
        state_var_NS = main_C_15;
      end
      main_C_15 : begin
        fsm_output = 8'b00010010;
        state_var_NS = main_C_16;
      end
      main_C_16 : begin
        fsm_output = 8'b00010011;
        state_var_NS = main_C_17;
      end
      main_C_17 : begin
        fsm_output = 8'b00010100;
        state_var_NS = main_C_18;
      end
      main_C_18 : begin
        fsm_output = 8'b00010101;
        state_var_NS = main_C_19;
      end
      main_C_19 : begin
        fsm_output = 8'b00010110;
        state_var_NS = main_C_20;
      end
      main_C_20 : begin
        fsm_output = 8'b00010111;
        state_var_NS = main_C_21;
      end
      main_C_21 : begin
        fsm_output = 8'b00011000;
        state_var_NS = main_C_22;
      end
      main_C_22 : begin
        fsm_output = 8'b00011001;
        state_var_NS = main_C_23;
      end
      main_C_23 : begin
        fsm_output = 8'b00011010;
        state_var_NS = main_C_24;
      end
      main_C_24 : begin
        fsm_output = 8'b00011011;
        state_var_NS = main_C_25;
      end
      main_C_25 : begin
        fsm_output = 8'b00011100;
        state_var_NS = main_C_26;
      end
      main_C_26 : begin
        fsm_output = 8'b00011101;
        state_var_NS = main_C_27;
      end
      main_C_27 : begin
        fsm_output = 8'b00011110;
        state_var_NS = main_C_28;
      end
      main_C_28 : begin
        fsm_output = 8'b00011111;
        state_var_NS = main_C_29;
      end
      main_C_29 : begin
        fsm_output = 8'b00100000;
        state_var_NS = main_C_30;
      end
      main_C_30 : begin
        fsm_output = 8'b00100001;
        state_var_NS = main_C_31;
      end
      main_C_31 : begin
        fsm_output = 8'b00100010;
        state_var_NS = main_C_32;
      end
      main_C_32 : begin
        fsm_output = 8'b00100011;
        state_var_NS = main_C_33;
      end
      main_C_33 : begin
        fsm_output = 8'b00100100;
        state_var_NS = main_C_34;
      end
      main_C_34 : begin
        fsm_output = 8'b00100101;
        state_var_NS = main_C_35;
      end
      main_C_35 : begin
        fsm_output = 8'b00100110;
        state_var_NS = main_C_36;
      end
      main_C_36 : begin
        fsm_output = 8'b00100111;
        state_var_NS = main_C_37;
      end
      main_C_37 : begin
        fsm_output = 8'b00101000;
        state_var_NS = main_C_38;
      end
      main_C_38 : begin
        fsm_output = 8'b00101001;
        state_var_NS = main_C_39;
      end
      main_C_39 : begin
        fsm_output = 8'b00101010;
        state_var_NS = main_C_40;
      end
      main_C_40 : begin
        fsm_output = 8'b00101011;
        state_var_NS = main_C_41;
      end
      main_C_41 : begin
        fsm_output = 8'b00101100;
        state_var_NS = main_C_42;
      end
      main_C_42 : begin
        fsm_output = 8'b00101101;
        state_var_NS = main_C_43;
      end
      main_C_43 : begin
        fsm_output = 8'b00101110;
        state_var_NS = main_C_44;
      end
      main_C_44 : begin
        fsm_output = 8'b00101111;
        state_var_NS = main_C_45;
      end
      main_C_45 : begin
        fsm_output = 8'b00110000;
        state_var_NS = main_C_46;
      end
      main_C_46 : begin
        fsm_output = 8'b00110001;
        state_var_NS = main_C_47;
      end
      main_C_47 : begin
        fsm_output = 8'b00110010;
        state_var_NS = main_C_48;
      end
      main_C_48 : begin
        fsm_output = 8'b00110011;
        state_var_NS = main_C_49;
      end
      main_C_49 : begin
        fsm_output = 8'b00110100;
        state_var_NS = main_C_50;
      end
      main_C_50 : begin
        fsm_output = 8'b00110101;
        state_var_NS = main_C_51;
      end
      main_C_51 : begin
        fsm_output = 8'b00110110;
        state_var_NS = main_C_52;
      end
      main_C_52 : begin
        fsm_output = 8'b00110111;
        state_var_NS = main_C_53;
      end
      main_C_53 : begin
        fsm_output = 8'b00111000;
        state_var_NS = main_C_54;
      end
      main_C_54 : begin
        fsm_output = 8'b00111001;
        state_var_NS = main_C_55;
      end
      main_C_55 : begin
        fsm_output = 8'b00111010;
        state_var_NS = main_C_56;
      end
      main_C_56 : begin
        fsm_output = 8'b00111011;
        state_var_NS = main_C_57;
      end
      main_C_57 : begin
        fsm_output = 8'b00111100;
        state_var_NS = main_C_58;
      end
      main_C_58 : begin
        fsm_output = 8'b00111101;
        state_var_NS = main_C_59;
      end
      main_C_59 : begin
        fsm_output = 8'b00111110;
        state_var_NS = main_C_60;
      end
      main_C_60 : begin
        fsm_output = 8'b00111111;
        state_var_NS = main_C_61;
      end
      main_C_61 : begin
        fsm_output = 8'b01000000;
        state_var_NS = main_C_62;
      end
      main_C_62 : begin
        fsm_output = 8'b01000001;
        state_var_NS = main_C_63;
      end
      main_C_63 : begin
        fsm_output = 8'b01000010;
        state_var_NS = main_C_64;
      end
      main_C_64 : begin
        fsm_output = 8'b01000011;
        state_var_NS = InitAccumLoop_1_C_0;
      end
      InitAccumLoop_1_C_0 : begin
        fsm_output = 8'b01000100;
        if ( InitAccumLoop_1_C_0_tr0 ) begin
          state_var_NS = ReuseLoop_1_C_0;
        end
        else begin
          state_var_NS = InitAccumLoop_1_C_0;
        end
      end
      ReuseLoop_1_C_0 : begin
        fsm_output = 8'b01000101;
        if ( ReuseLoop_1_C_0_tr0 ) begin
          state_var_NS = main_C_65;
        end
        else begin
          state_var_NS = ReuseLoop_1_C_0;
        end
      end
      main_C_65 : begin
        fsm_output = 8'b01000110;
        state_var_NS = main_C_66;
      end
      main_C_66 : begin
        fsm_output = 8'b01000111;
        state_var_NS = main_C_67;
      end
      main_C_67 : begin
        fsm_output = 8'b01001000;
        state_var_NS = main_C_68;
      end
      main_C_68 : begin
        fsm_output = 8'b01001001;
        state_var_NS = main_C_69;
      end
      main_C_69 : begin
        fsm_output = 8'b01001010;
        state_var_NS = main_C_70;
      end
      main_C_70 : begin
        fsm_output = 8'b01001011;
        state_var_NS = main_C_71;
      end
      main_C_71 : begin
        fsm_output = 8'b01001100;
        state_var_NS = main_C_72;
      end
      main_C_72 : begin
        fsm_output = 8'b01001101;
        state_var_NS = main_C_73;
      end
      main_C_73 : begin
        fsm_output = 8'b01001110;
        state_var_NS = main_C_74;
      end
      main_C_74 : begin
        fsm_output = 8'b01001111;
        state_var_NS = main_C_75;
      end
      main_C_75 : begin
        fsm_output = 8'b01010000;
        state_var_NS = main_C_76;
      end
      main_C_76 : begin
        fsm_output = 8'b01010001;
        state_var_NS = main_C_77;
      end
      main_C_77 : begin
        fsm_output = 8'b01010010;
        state_var_NS = main_C_78;
      end
      main_C_78 : begin
        fsm_output = 8'b01010011;
        state_var_NS = main_C_79;
      end
      main_C_79 : begin
        fsm_output = 8'b01010100;
        state_var_NS = main_C_80;
      end
      main_C_80 : begin
        fsm_output = 8'b01010101;
        state_var_NS = main_C_81;
      end
      main_C_81 : begin
        fsm_output = 8'b01010110;
        state_var_NS = main_C_82;
      end
      main_C_82 : begin
        fsm_output = 8'b01010111;
        state_var_NS = main_C_83;
      end
      main_C_83 : begin
        fsm_output = 8'b01011000;
        state_var_NS = main_C_84;
      end
      main_C_84 : begin
        fsm_output = 8'b01011001;
        state_var_NS = main_C_85;
      end
      main_C_85 : begin
        fsm_output = 8'b01011010;
        state_var_NS = main_C_86;
      end
      main_C_86 : begin
        fsm_output = 8'b01011011;
        state_var_NS = main_C_87;
      end
      main_C_87 : begin
        fsm_output = 8'b01011100;
        state_var_NS = main_C_88;
      end
      main_C_88 : begin
        fsm_output = 8'b01011101;
        state_var_NS = main_C_89;
      end
      main_C_89 : begin
        fsm_output = 8'b01011110;
        state_var_NS = main_C_90;
      end
      main_C_90 : begin
        fsm_output = 8'b01011111;
        state_var_NS = main_C_91;
      end
      main_C_91 : begin
        fsm_output = 8'b01100000;
        state_var_NS = main_C_92;
      end
      main_C_92 : begin
        fsm_output = 8'b01100001;
        state_var_NS = main_C_93;
      end
      main_C_93 : begin
        fsm_output = 8'b01100010;
        state_var_NS = main_C_94;
      end
      main_C_94 : begin
        fsm_output = 8'b01100011;
        state_var_NS = main_C_95;
      end
      main_C_95 : begin
        fsm_output = 8'b01100100;
        state_var_NS = main_C_96;
      end
      main_C_96 : begin
        fsm_output = 8'b01100101;
        state_var_NS = main_C_97;
      end
      main_C_97 : begin
        fsm_output = 8'b01100110;
        state_var_NS = main_C_98;
      end
      main_C_98 : begin
        fsm_output = 8'b01100111;
        state_var_NS = main_C_99;
      end
      main_C_99 : begin
        fsm_output = 8'b01101000;
        state_var_NS = main_C_100;
      end
      main_C_100 : begin
        fsm_output = 8'b01101001;
        state_var_NS = main_C_101;
      end
      main_C_101 : begin
        fsm_output = 8'b01101010;
        state_var_NS = main_C_102;
      end
      main_C_102 : begin
        fsm_output = 8'b01101011;
        state_var_NS = main_C_103;
      end
      main_C_103 : begin
        fsm_output = 8'b01101100;
        state_var_NS = main_C_104;
      end
      main_C_104 : begin
        fsm_output = 8'b01101101;
        state_var_NS = main_C_105;
      end
      main_C_105 : begin
        fsm_output = 8'b01101110;
        state_var_NS = main_C_106;
      end
      main_C_106 : begin
        fsm_output = 8'b01101111;
        state_var_NS = main_C_107;
      end
      main_C_107 : begin
        fsm_output = 8'b01110000;
        state_var_NS = main_C_108;
      end
      main_C_108 : begin
        fsm_output = 8'b01110001;
        state_var_NS = main_C_109;
      end
      main_C_109 : begin
        fsm_output = 8'b01110010;
        state_var_NS = main_C_110;
      end
      main_C_110 : begin
        fsm_output = 8'b01110011;
        state_var_NS = main_C_111;
      end
      main_C_111 : begin
        fsm_output = 8'b01110100;
        state_var_NS = main_C_112;
      end
      main_C_112 : begin
        fsm_output = 8'b01110101;
        state_var_NS = main_C_113;
      end
      main_C_113 : begin
        fsm_output = 8'b01110110;
        state_var_NS = main_C_114;
      end
      main_C_114 : begin
        fsm_output = 8'b01110111;
        state_var_NS = main_C_115;
      end
      main_C_115 : begin
        fsm_output = 8'b01111000;
        state_var_NS = main_C_116;
      end
      main_C_116 : begin
        fsm_output = 8'b01111001;
        state_var_NS = main_C_117;
      end
      main_C_117 : begin
        fsm_output = 8'b01111010;
        state_var_NS = main_C_118;
      end
      main_C_118 : begin
        fsm_output = 8'b01111011;
        state_var_NS = main_C_119;
      end
      main_C_119 : begin
        fsm_output = 8'b01111100;
        state_var_NS = main_C_120;
      end
      main_C_120 : begin
        fsm_output = 8'b01111101;
        state_var_NS = main_C_121;
      end
      main_C_121 : begin
        fsm_output = 8'b01111110;
        state_var_NS = main_C_122;
      end
      main_C_122 : begin
        fsm_output = 8'b01111111;
        state_var_NS = main_C_123;
      end
      main_C_123 : begin
        fsm_output = 8'b10000000;
        state_var_NS = main_C_124;
      end
      main_C_124 : begin
        fsm_output = 8'b10000001;
        state_var_NS = main_C_125;
      end
      main_C_125 : begin
        fsm_output = 8'b10000010;
        state_var_NS = main_C_126;
      end
      main_C_126 : begin
        fsm_output = 8'b10000011;
        state_var_NS = main_C_127;
      end
      main_C_127 : begin
        fsm_output = 8'b10000100;
        state_var_NS = main_C_128;
      end
      main_C_128 : begin
        fsm_output = 8'b10000101;
        state_var_NS = InitAccumLoop_2_C_0;
      end
      InitAccumLoop_2_C_0 : begin
        fsm_output = 8'b10000110;
        if ( InitAccumLoop_2_C_0_tr0 ) begin
          state_var_NS = ReuseLoop_2_C_0;
        end
        else begin
          state_var_NS = InitAccumLoop_2_C_0;
        end
      end
      ReuseLoop_2_C_0 : begin
        fsm_output = 8'b10000111;
        if ( ReuseLoop_2_C_0_tr0 ) begin
          state_var_NS = main_C_129;
        end
        else begin
          state_var_NS = ReuseLoop_2_C_0;
        end
      end
      main_C_129 : begin
        fsm_output = 8'b10001000;
        state_var_NS = main_C_130;
      end
      main_C_130 : begin
        fsm_output = 8'b10001001;
        state_var_NS = main_C_131;
      end
      main_C_131 : begin
        fsm_output = 8'b10001010;
        state_var_NS = main_C_132;
      end
      main_C_132 : begin
        fsm_output = 8'b10001011;
        state_var_NS = main_C_133;
      end
      main_C_133 : begin
        fsm_output = 8'b10001100;
        state_var_NS = main_C_134;
      end
      main_C_134 : begin
        fsm_output = 8'b10001101;
        state_var_NS = main_C_135;
      end
      main_C_135 : begin
        fsm_output = 8'b10001110;
        state_var_NS = main_C_136;
      end
      main_C_136 : begin
        fsm_output = 8'b10001111;
        state_var_NS = main_C_137;
      end
      main_C_137 : begin
        fsm_output = 8'b10010000;
        state_var_NS = main_C_138;
      end
      main_C_138 : begin
        fsm_output = 8'b10010001;
        state_var_NS = main_C_139;
      end
      main_C_139 : begin
        fsm_output = 8'b10010010;
        state_var_NS = main_C_140;
      end
      main_C_140 : begin
        fsm_output = 8'b10010011;
        state_var_NS = main_C_141;
      end
      main_C_141 : begin
        fsm_output = 8'b10010100;
        state_var_NS = main_C_142;
      end
      main_C_142 : begin
        fsm_output = 8'b10010101;
        state_var_NS = main_C_143;
      end
      main_C_143 : begin
        fsm_output = 8'b10010110;
        state_var_NS = main_C_144;
      end
      main_C_144 : begin
        fsm_output = 8'b10010111;
        state_var_NS = main_C_145;
      end
      main_C_145 : begin
        fsm_output = 8'b10011000;
        state_var_NS = main_C_146;
      end
      main_C_146 : begin
        fsm_output = 8'b10011001;
        state_var_NS = main_C_147;
      end
      main_C_147 : begin
        fsm_output = 8'b10011010;
        state_var_NS = main_C_148;
      end
      main_C_148 : begin
        fsm_output = 8'b10011011;
        state_var_NS = main_C_149;
      end
      main_C_149 : begin
        fsm_output = 8'b10011100;
        state_var_NS = main_C_150;
      end
      main_C_150 : begin
        fsm_output = 8'b10011101;
        state_var_NS = nnet_softmax_layer6_t_result_t_softmax_config7_for_1_C_0;
      end
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_C_0 : begin
        fsm_output = 8'b10011110;
        if ( nnet_softmax_layer6_t_result_t_softmax_config7_for_1_C_0_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = nnet_softmax_layer6_t_result_t_softmax_config7_for_1_C_0;
        end
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 8'b00000000;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_staller
// ------------------------------------------------------------------


module mnist_mlp_core_staller (
  clk, rst, core_wen, core_wten, input1_rsci_wen_comp, layer7_out_rsci_wen_comp,
      const_size_in_1_rsci_wen_comp, const_size_out_1_rsci_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  input input1_rsci_wen_comp;
  input layer7_out_rsci_wen_comp;
  input const_size_in_1_rsci_wen_comp;
  input const_size_out_1_rsci_wen_comp;


  // Interconnect Declarations
  reg core_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign core_wen = input1_rsci_wen_comp & layer7_out_rsci_wen_comp & const_size_in_1_rsci_wen_comp
      & const_size_out_1_rsci_wen_comp;
  assign core_wten = core_wten_reg;
  always @(posedge clk) begin
    if ( rst ) begin
      core_wten_reg <= 1'b0;
    end
    else begin
      core_wten_reg <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_w6_rsci_1_w6_rsc_wait_dp
// ------------------------------------------------------------------


module mnist_mlp_core_w6_rsci_1_w6_rsc_wait_dp (
  clk, rst, w6_rsci_adra_d, w6_rsci_qa_d, w6_rsci_qa_d_mxwt, w6_rsci_biwt, w6_rsci_bdwt,
      w6_rsci_adra_d_core_sct, w6_rsci_adra_d_core_pff
);
  input clk;
  input rst;
  output [19:0] w6_rsci_adra_d;
  input [35:0] w6_rsci_qa_d;
  output [35:0] w6_rsci_qa_d_mxwt;
  input w6_rsci_biwt;
  input w6_rsci_bdwt;
  input [1:0] w6_rsci_adra_d_core_sct;
  input [19:0] w6_rsci_adra_d_core_pff;


  // Interconnect Declarations
  reg w6_rsci_bcwt;
  reg w6_rsci_bcwt_1;
  reg [17:0] w6_rsci_qa_d_bfwt_35_18;
  reg [17:0] w6_rsci_qa_d_bfwt_17_0;

  wire[17:0] MultLoop_2_mux_nl;
  wire[17:0] MultLoop_2_mux_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign MultLoop_2_mux_nl = MUX_v_18_2_2((w6_rsci_qa_d[35:18]), w6_rsci_qa_d_bfwt_35_18,
      w6_rsci_bcwt_1);
  assign MultLoop_2_mux_1_nl = MUX_v_18_2_2((w6_rsci_qa_d[17:0]), w6_rsci_qa_d_bfwt_17_0,
      w6_rsci_bcwt);
  assign w6_rsci_qa_d_mxwt = {(MultLoop_2_mux_nl) , (MultLoop_2_mux_1_nl)};
  assign w6_rsci_adra_d = {(w6_rsci_adra_d_core_pff[19:10]) , (~ (w6_rsci_adra_d_core_sct[0]))
      , (w6_rsci_adra_d_core_pff[8:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      w6_rsci_bcwt <= 1'b0;
      w6_rsci_bcwt_1 <= 1'b0;
    end
    else begin
      w6_rsci_bcwt <= ~((~(w6_rsci_bcwt | w6_rsci_biwt)) | w6_rsci_bdwt);
      w6_rsci_bcwt_1 <= ~((~(w6_rsci_bcwt_1 | w6_rsci_biwt)) | w6_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      w6_rsci_qa_d_bfwt_35_18 <= 18'b000000000000000000;
    end
    else if ( ~ w6_rsci_bcwt_1 ) begin
      w6_rsci_qa_d_bfwt_35_18 <= w6_rsci_qa_d_mxwt[35:18];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      w6_rsci_qa_d_bfwt_17_0 <= 18'b000000000000000000;
    end
    else if ( ~ w6_rsci_bcwt ) begin
      w6_rsci_qa_d_bfwt_17_0 <= w6_rsci_qa_d_mxwt[17:0];
    end
  end

  function automatic [17:0] MUX_v_18_2_2;
    input [17:0] input_0;
    input [17:0] input_1;
    input [0:0] sel;
    reg [17:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_18_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_w6_rsci_1_w6_rsc_wait_ctrl
// ------------------------------------------------------------------


module mnist_mlp_core_w6_rsci_1_w6_rsc_wait_ctrl (
  core_wen, core_wten, w6_rsci_oswt, w6_rsci_adra_d_core_psct, w6_rsci_ena_d_core_psct,
      w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct, w6_rsci_biwt, w6_rsci_bdwt,
      w6_rsci_adra_d_core_sct, w6_rsci_ena_d_core_sct, w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      w6_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input w6_rsci_oswt;
  input [1:0] w6_rsci_adra_d_core_psct;
  input [1:0] w6_rsci_ena_d_core_psct;
  input [1:0] w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  output w6_rsci_biwt;
  output w6_rsci_bdwt;
  output [1:0] w6_rsci_adra_d_core_sct;
  output [1:0] w6_rsci_ena_d_core_sct;
  output [1:0] w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  input w6_rsci_oswt_pff;


  // Interconnect Declarations
  wire w6_rsci_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign w6_rsci_bdwt = w6_rsci_oswt & core_wen;
  assign w6_rsci_biwt = (~ core_wten) & w6_rsci_oswt;
  assign w6_rsci_adra_d_core_sct = w6_rsci_adra_d_core_psct & ({w6_rsci_dswt_pff
      , w6_rsci_dswt_pff});
  assign w6_rsci_dswt_pff = core_wen & w6_rsci_oswt_pff;
  assign w6_rsci_ena_d_core_sct = w6_rsci_ena_d_core_psct & ({w6_rsci_dswt_pff ,
      w6_rsci_dswt_pff});
  assign w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & ({w6_rsci_dswt_pff , w6_rsci_dswt_pff});
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_w4_rsci_1_w4_rsc_wait_dp
// ------------------------------------------------------------------


module mnist_mlp_core_w4_rsci_1_w4_rsc_wait_dp (
  clk, rst, w4_rsci_adra_d, w4_rsci_qa_d, w4_rsci_qa_d_mxwt, w4_rsci_biwt, w4_rsci_bdwt,
      w4_rsci_adra_d_core_sct_pff, w4_rsci_adra_d_core_pff
);
  input clk;
  input rst;
  output [23:0] w4_rsci_adra_d;
  input [35:0] w4_rsci_qa_d;
  output [35:0] w4_rsci_qa_d_mxwt;
  input w4_rsci_biwt;
  input w4_rsci_bdwt;
  input [1:0] w4_rsci_adra_d_core_sct_pff;
  input [23:0] w4_rsci_adra_d_core_pff;


  // Interconnect Declarations
  reg w4_rsci_bcwt;
  reg w4_rsci_bcwt_1;
  reg [17:0] w4_rsci_qa_d_bfwt_35_18;
  reg [17:0] w4_rsci_qa_d_bfwt_17_0;

  wire[17:0] MultLoop_1_mux_nl;
  wire[17:0] MultLoop_1_mux_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign MultLoop_1_mux_nl = MUX_v_18_2_2((w4_rsci_qa_d[35:18]), w4_rsci_qa_d_bfwt_35_18,
      w4_rsci_bcwt_1);
  assign MultLoop_1_mux_1_nl = MUX_v_18_2_2((w4_rsci_qa_d[17:0]), w4_rsci_qa_d_bfwt_17_0,
      w4_rsci_bcwt);
  assign w4_rsci_qa_d_mxwt = {(MultLoop_1_mux_nl) , (MultLoop_1_mux_1_nl)};
  assign w4_rsci_adra_d = {(w4_rsci_adra_d_core_sct_pff[1]) , (w4_rsci_adra_d_core_pff[22:12])
      , (~ (w4_rsci_adra_d_core_sct_pff[0])) , (w4_rsci_adra_d_core_pff[10:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      w4_rsci_bcwt <= 1'b0;
      w4_rsci_bcwt_1 <= 1'b0;
    end
    else begin
      w4_rsci_bcwt <= ~((~(w4_rsci_bcwt | w4_rsci_biwt)) | w4_rsci_bdwt);
      w4_rsci_bcwt_1 <= ~((~(w4_rsci_bcwt_1 | w4_rsci_biwt)) | w4_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      w4_rsci_qa_d_bfwt_35_18 <= 18'b000000000000000000;
    end
    else if ( ~ w4_rsci_bcwt_1 ) begin
      w4_rsci_qa_d_bfwt_35_18 <= w4_rsci_qa_d_mxwt[35:18];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      w4_rsci_qa_d_bfwt_17_0 <= 18'b000000000000000000;
    end
    else if ( ~ w4_rsci_bcwt ) begin
      w4_rsci_qa_d_bfwt_17_0 <= w4_rsci_qa_d_mxwt[17:0];
    end
  end

  function automatic [17:0] MUX_v_18_2_2;
    input [17:0] input_0;
    input [17:0] input_1;
    input [0:0] sel;
    reg [17:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_18_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_w4_rsci_1_w4_rsc_wait_ctrl
// ------------------------------------------------------------------


module mnist_mlp_core_w4_rsci_1_w4_rsc_wait_ctrl (
  core_wen, core_wten, w4_rsci_oswt, w4_rsci_ena_d_core_psct, w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      w4_rsci_biwt, w4_rsci_bdwt, w4_rsci_ena_d_core_sct, w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      w4_rsci_adra_d_core_sct_pff, w4_rsci_adra_d_core_psct_pff, w4_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input w4_rsci_oswt;
  input [1:0] w4_rsci_ena_d_core_psct;
  input [1:0] w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  output w4_rsci_biwt;
  output w4_rsci_bdwt;
  output [1:0] w4_rsci_ena_d_core_sct;
  output [1:0] w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output [1:0] w4_rsci_adra_d_core_sct_pff;
  input [1:0] w4_rsci_adra_d_core_psct_pff;
  input w4_rsci_oswt_pff;


  // Interconnect Declarations
  wire w4_rsci_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign w4_rsci_bdwt = w4_rsci_oswt & core_wen;
  assign w4_rsci_biwt = (~ core_wten) & w4_rsci_oswt;
  assign w4_rsci_adra_d_core_sct_pff = w4_rsci_adra_d_core_psct_pff & ({w4_rsci_dswt_pff
      , w4_rsci_dswt_pff});
  assign w4_rsci_dswt_pff = core_wen & w4_rsci_oswt_pff;
  assign w4_rsci_ena_d_core_sct = w4_rsci_ena_d_core_psct & ({w4_rsci_dswt_pff ,
      w4_rsci_dswt_pff});
  assign w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & ({w4_rsci_dswt_pff , w4_rsci_dswt_pff});
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_w2_rsci_1_w2_rsc_wait_dp
// ------------------------------------------------------------------


module mnist_mlp_core_w2_rsci_1_w2_rsc_wait_dp (
  clk, rst, w2_rsci_adra_d, w2_rsci_qa_d, w2_rsci_qa_d_mxwt, w2_rsci_biwt, w2_rsci_bdwt,
      w2_rsci_adra_d_core_sct, w2_rsci_adra_d_core_pff
);
  input clk;
  input rst;
  output [31:0] w2_rsci_adra_d;
  input [35:0] w2_rsci_qa_d;
  output [35:0] w2_rsci_qa_d_mxwt;
  input w2_rsci_biwt;
  input w2_rsci_bdwt;
  input [1:0] w2_rsci_adra_d_core_sct;
  input [31:0] w2_rsci_adra_d_core_pff;


  // Interconnect Declarations
  reg w2_rsci_bcwt;
  reg w2_rsci_bcwt_1;
  reg [17:0] w2_rsci_qa_d_bfwt_35_18;
  reg [17:0] w2_rsci_qa_d_bfwt_17_0;

  wire[17:0] MultLoop_mux_1_nl;
  wire[17:0] MultLoop_mux_2_nl;

  // Interconnect Declarations for Component Instantiations 
  assign MultLoop_mux_1_nl = MUX_v_18_2_2((w2_rsci_qa_d[35:18]), w2_rsci_qa_d_bfwt_35_18,
      w2_rsci_bcwt_1);
  assign MultLoop_mux_2_nl = MUX_v_18_2_2((w2_rsci_qa_d[17:0]), w2_rsci_qa_d_bfwt_17_0,
      w2_rsci_bcwt);
  assign w2_rsci_qa_d_mxwt = {(MultLoop_mux_1_nl) , (MultLoop_mux_2_nl)};
  assign w2_rsci_adra_d = {(w2_rsci_adra_d_core_pff[31:16]) , (~ (w2_rsci_adra_d_core_sct[0]))
      , (w2_rsci_adra_d_core_pff[14:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      w2_rsci_bcwt <= 1'b0;
      w2_rsci_bcwt_1 <= 1'b0;
    end
    else begin
      w2_rsci_bcwt <= ~((~(w2_rsci_bcwt | w2_rsci_biwt)) | w2_rsci_bdwt);
      w2_rsci_bcwt_1 <= ~((~(w2_rsci_bcwt_1 | w2_rsci_biwt)) | w2_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      w2_rsci_qa_d_bfwt_35_18 <= 18'b000000000000000000;
    end
    else if ( ~ w2_rsci_bcwt_1 ) begin
      w2_rsci_qa_d_bfwt_35_18 <= w2_rsci_qa_d_mxwt[35:18];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      w2_rsci_qa_d_bfwt_17_0 <= 18'b000000000000000000;
    end
    else if ( ~ w2_rsci_bcwt ) begin
      w2_rsci_qa_d_bfwt_17_0 <= w2_rsci_qa_d_mxwt[17:0];
    end
  end

  function automatic [17:0] MUX_v_18_2_2;
    input [17:0] input_0;
    input [17:0] input_1;
    input [0:0] sel;
    reg [17:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_18_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_w2_rsci_1_w2_rsc_wait_ctrl
// ------------------------------------------------------------------


module mnist_mlp_core_w2_rsci_1_w2_rsc_wait_ctrl (
  core_wen, core_wten, w2_rsci_oswt, w2_rsci_adra_d_core_psct, w2_rsci_ena_d_core_psct,
      w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct, w2_rsci_biwt, w2_rsci_bdwt,
      w2_rsci_adra_d_core_sct, w2_rsci_ena_d_core_sct, w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      w2_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input w2_rsci_oswt;
  input [1:0] w2_rsci_adra_d_core_psct;
  input [1:0] w2_rsci_ena_d_core_psct;
  input [1:0] w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  output w2_rsci_biwt;
  output w2_rsci_bdwt;
  output [1:0] w2_rsci_adra_d_core_sct;
  output [1:0] w2_rsci_ena_d_core_sct;
  output [1:0] w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  input w2_rsci_oswt_pff;


  // Interconnect Declarations
  wire w2_rsci_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign w2_rsci_bdwt = w2_rsci_oswt & core_wen;
  assign w2_rsci_biwt = (~ core_wten) & w2_rsci_oswt;
  assign w2_rsci_adra_d_core_sct = w2_rsci_adra_d_core_psct & ({w2_rsci_dswt_pff
      , w2_rsci_dswt_pff});
  assign w2_rsci_dswt_pff = core_wen & w2_rsci_oswt_pff;
  assign w2_rsci_ena_d_core_sct = w2_rsci_ena_d_core_psct & ({w2_rsci_dswt_pff ,
      w2_rsci_dswt_pff});
  assign w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & ({w2_rsci_dswt_pff , w2_rsci_dswt_pff});
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_dp
// ------------------------------------------------------------------


module mnist_mlp_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_dp (
  clk, rst, const_size_out_1_rsci_oswt, const_size_out_1_rsci_wen_comp, const_size_out_1_rsci_biwt,
      const_size_out_1_rsci_bdwt, const_size_out_1_rsci_bcwt
);
  input clk;
  input rst;
  input const_size_out_1_rsci_oswt;
  output const_size_out_1_rsci_wen_comp;
  input const_size_out_1_rsci_biwt;
  input const_size_out_1_rsci_bdwt;
  output const_size_out_1_rsci_bcwt;
  reg const_size_out_1_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_out_1_rsci_wen_comp = (~ const_size_out_1_rsci_oswt) | const_size_out_1_rsci_biwt
      | const_size_out_1_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      const_size_out_1_rsci_bcwt <= 1'b0;
    end
    else begin
      const_size_out_1_rsci_bcwt <= ~((~(const_size_out_1_rsci_bcwt | const_size_out_1_rsci_biwt))
          | const_size_out_1_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module mnist_mlp_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl (
  core_wen, const_size_out_1_rsci_oswt, const_size_out_1_rsci_irdy, const_size_out_1_rsci_biwt,
      const_size_out_1_rsci_bdwt, const_size_out_1_rsci_bcwt, const_size_out_1_rsci_ivld_core_sct
);
  input core_wen;
  input const_size_out_1_rsci_oswt;
  input const_size_out_1_rsci_irdy;
  output const_size_out_1_rsci_biwt;
  output const_size_out_1_rsci_bdwt;
  input const_size_out_1_rsci_bcwt;
  output const_size_out_1_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire const_size_out_1_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign const_size_out_1_rsci_bdwt = const_size_out_1_rsci_oswt & core_wen;
  assign const_size_out_1_rsci_biwt = const_size_out_1_rsci_ogwt & const_size_out_1_rsci_irdy;
  assign const_size_out_1_rsci_ogwt = const_size_out_1_rsci_oswt & (~ const_size_out_1_rsci_bcwt);
  assign const_size_out_1_rsci_ivld_core_sct = const_size_out_1_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_dp
// ------------------------------------------------------------------


module mnist_mlp_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_dp (
  clk, rst, const_size_in_1_rsci_oswt, const_size_in_1_rsci_wen_comp, const_size_in_1_rsci_biwt,
      const_size_in_1_rsci_bdwt, const_size_in_1_rsci_bcwt
);
  input clk;
  input rst;
  input const_size_in_1_rsci_oswt;
  output const_size_in_1_rsci_wen_comp;
  input const_size_in_1_rsci_biwt;
  input const_size_in_1_rsci_bdwt;
  output const_size_in_1_rsci_bcwt;
  reg const_size_in_1_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_in_1_rsci_wen_comp = (~ const_size_in_1_rsci_oswt) | const_size_in_1_rsci_biwt
      | const_size_in_1_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      const_size_in_1_rsci_bcwt <= 1'b0;
    end
    else begin
      const_size_in_1_rsci_bcwt <= ~((~(const_size_in_1_rsci_bcwt | const_size_in_1_rsci_biwt))
          | const_size_in_1_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module mnist_mlp_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl (
  core_wen, const_size_in_1_rsci_oswt, const_size_in_1_rsci_irdy, const_size_in_1_rsci_biwt,
      const_size_in_1_rsci_bdwt, const_size_in_1_rsci_bcwt, const_size_in_1_rsci_ivld_core_sct
);
  input core_wen;
  input const_size_in_1_rsci_oswt;
  input const_size_in_1_rsci_irdy;
  output const_size_in_1_rsci_biwt;
  output const_size_in_1_rsci_bdwt;
  input const_size_in_1_rsci_bcwt;
  output const_size_in_1_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire const_size_in_1_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign const_size_in_1_rsci_bdwt = const_size_in_1_rsci_oswt & core_wen;
  assign const_size_in_1_rsci_biwt = const_size_in_1_rsci_ogwt & const_size_in_1_rsci_irdy;
  assign const_size_in_1_rsci_ogwt = const_size_in_1_rsci_oswt & (~ const_size_in_1_rsci_bcwt);
  assign const_size_in_1_rsci_ivld_core_sct = const_size_in_1_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_layer7_out_rsci_layer7_out_rsc_wait_dp
// ------------------------------------------------------------------


module mnist_mlp_core_layer7_out_rsci_layer7_out_rsc_wait_dp (
  clk, rst, layer7_out_rsci_oswt, layer7_out_rsci_wen_comp, layer7_out_rsci_biwt,
      layer7_out_rsci_bdwt, layer7_out_rsci_bcwt
);
  input clk;
  input rst;
  input layer7_out_rsci_oswt;
  output layer7_out_rsci_wen_comp;
  input layer7_out_rsci_biwt;
  input layer7_out_rsci_bdwt;
  output layer7_out_rsci_bcwt;
  reg layer7_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign layer7_out_rsci_wen_comp = (~ layer7_out_rsci_oswt) | layer7_out_rsci_biwt
      | layer7_out_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      layer7_out_rsci_bcwt <= 1'b0;
    end
    else begin
      layer7_out_rsci_bcwt <= ~((~(layer7_out_rsci_bcwt | layer7_out_rsci_biwt))
          | layer7_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_layer7_out_rsci_layer7_out_rsc_wait_ctrl
// ------------------------------------------------------------------


module mnist_mlp_core_layer7_out_rsci_layer7_out_rsc_wait_ctrl (
  core_wen, layer7_out_rsci_oswt, layer7_out_rsci_irdy, layer7_out_rsci_biwt, layer7_out_rsci_bdwt,
      layer7_out_rsci_bcwt, layer7_out_rsci_ivld_core_sct
);
  input core_wen;
  input layer7_out_rsci_oswt;
  input layer7_out_rsci_irdy;
  output layer7_out_rsci_biwt;
  output layer7_out_rsci_bdwt;
  input layer7_out_rsci_bcwt;
  output layer7_out_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire layer7_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign layer7_out_rsci_bdwt = layer7_out_rsci_oswt & core_wen;
  assign layer7_out_rsci_biwt = layer7_out_rsci_ogwt & layer7_out_rsci_irdy;
  assign layer7_out_rsci_ogwt = layer7_out_rsci_oswt & (~ layer7_out_rsci_bcwt);
  assign layer7_out_rsci_ivld_core_sct = layer7_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_input1_rsci_input1_rsc_wait_dp
// ------------------------------------------------------------------


module mnist_mlp_core_input1_rsci_input1_rsc_wait_dp (
  clk, rst, input1_rsci_oswt, input1_rsci_wen_comp, input1_rsci_idat_mxwt, input1_rsci_biwt,
      input1_rsci_bdwt, input1_rsci_bcwt, input1_rsci_idat
);
  input clk;
  input rst;
  input input1_rsci_oswt;
  output input1_rsci_wen_comp;
  output [14111:0] input1_rsci_idat_mxwt;
  input input1_rsci_biwt;
  input input1_rsci_bdwt;
  output input1_rsci_bcwt;
  reg input1_rsci_bcwt;
  input [14111:0] input1_rsci_idat;


  // Interconnect Declarations
  reg [14111:0] input1_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign input1_rsci_wen_comp = (~ input1_rsci_oswt) | input1_rsci_biwt | input1_rsci_bcwt;
  assign input1_rsci_idat_mxwt = MUX_v_14112_2_2(input1_rsci_idat, input1_rsci_idat_bfwt,
      input1_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      input1_rsci_bcwt <= 1'b0;
    end
    else begin
      input1_rsci_bcwt <= ~((~(input1_rsci_bcwt | input1_rsci_biwt)) | input1_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      input1_rsci_idat_bfwt <= {882'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 882'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 882'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 882'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 882'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 882'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 882'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 882'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 882'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 882'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 882'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 882'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 882'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 882'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 882'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 882'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
    end
    else if ( ~ input1_rsci_bcwt ) begin
      input1_rsci_idat_bfwt <= input1_rsci_idat_mxwt;
    end
  end

  function automatic [14111:0] MUX_v_14112_2_2;
    input [14111:0] input_0;
    input [14111:0] input_1;
    input [0:0] sel;
    reg [14111:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14112_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_input1_rsci_input1_rsc_wait_ctrl
// ------------------------------------------------------------------


module mnist_mlp_core_input1_rsci_input1_rsc_wait_ctrl (
  core_wen, input1_rsci_oswt, input1_rsci_biwt, input1_rsci_bdwt, input1_rsci_bcwt,
      input1_rsci_irdy_core_sct, input1_rsci_ivld
);
  input core_wen;
  input input1_rsci_oswt;
  output input1_rsci_biwt;
  output input1_rsci_bdwt;
  input input1_rsci_bcwt;
  output input1_rsci_irdy_core_sct;
  input input1_rsci_ivld;


  // Interconnect Declarations
  wire input1_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign input1_rsci_bdwt = input1_rsci_oswt & core_wen;
  assign input1_rsci_biwt = input1_rsci_ogwt & input1_rsci_ivld;
  assign input1_rsci_ogwt = input1_rsci_oswt & (~ input1_rsci_bcwt);
  assign input1_rsci_irdy_core_sct = input1_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_w6_rsci_1
// ------------------------------------------------------------------


module mnist_mlp_core_w6_rsci_1 (
  clk, rst, w6_rsci_adra_d, w6_rsci_ena_d, w6_rsci_qa_d, w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, w6_rsci_oswt, w6_rsci_adra_d_core_psct, w6_rsci_ena_d_core_psct,
      w6_rsci_qa_d_mxwt, w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct, w6_rsci_adra_d_core_pff,
      w6_rsci_oswt_pff
);
  input clk;
  input rst;
  output [19:0] w6_rsci_adra_d;
  output [1:0] w6_rsci_ena_d;
  input [35:0] w6_rsci_qa_d;
  output [1:0] w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input w6_rsci_oswt;
  input [1:0] w6_rsci_adra_d_core_psct;
  input [1:0] w6_rsci_ena_d_core_psct;
  output [35:0] w6_rsci_qa_d_mxwt;
  input [1:0] w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input [19:0] w6_rsci_adra_d_core_pff;
  input w6_rsci_oswt_pff;


  // Interconnect Declarations
  wire w6_rsci_biwt;
  wire w6_rsci_bdwt;
  wire [1:0] w6_rsci_adra_d_core_sct;
  wire [1:0] w6_rsci_ena_d_core_sct;
  wire [1:0] w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire [19:0] w6_rsci_adra_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [19:0] nl_mnist_mlp_core_w6_rsci_1_w6_rsc_wait_dp_inst_w6_rsci_adra_d_core_pff;
  assign nl_mnist_mlp_core_w6_rsci_1_w6_rsc_wait_dp_inst_w6_rsci_adra_d_core_pff
      = {(w6_rsci_adra_d_core_pff[19:10]) , 1'b0 , (w6_rsci_adra_d_core_pff[8:0])};
  mnist_mlp_core_w6_rsci_1_w6_rsc_wait_ctrl mnist_mlp_core_w6_rsci_1_w6_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .w6_rsci_oswt(w6_rsci_oswt),
      .w6_rsci_adra_d_core_psct(w6_rsci_adra_d_core_psct),
      .w6_rsci_ena_d_core_psct(w6_rsci_ena_d_core_psct),
      .w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .w6_rsci_biwt(w6_rsci_biwt),
      .w6_rsci_bdwt(w6_rsci_bdwt),
      .w6_rsci_adra_d_core_sct(w6_rsci_adra_d_core_sct),
      .w6_rsci_ena_d_core_sct(w6_rsci_ena_d_core_sct),
      .w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .w6_rsci_oswt_pff(w6_rsci_oswt_pff)
    );
  mnist_mlp_core_w6_rsci_1_w6_rsc_wait_dp mnist_mlp_core_w6_rsci_1_w6_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .w6_rsci_adra_d(w6_rsci_adra_d_reg),
      .w6_rsci_qa_d(w6_rsci_qa_d),
      .w6_rsci_qa_d_mxwt(w6_rsci_qa_d_mxwt),
      .w6_rsci_biwt(w6_rsci_biwt),
      .w6_rsci_bdwt(w6_rsci_bdwt),
      .w6_rsci_adra_d_core_sct(w6_rsci_adra_d_core_sct),
      .w6_rsci_adra_d_core_pff(nl_mnist_mlp_core_w6_rsci_1_w6_rsc_wait_dp_inst_w6_rsci_adra_d_core_pff[19:0])
    );
  assign w6_rsci_adra_d = w6_rsci_adra_d_reg;
  assign w6_rsci_ena_d = w6_rsci_ena_d_core_sct;
  assign w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_w4_rsci_1
// ------------------------------------------------------------------


module mnist_mlp_core_w4_rsci_1 (
  clk, rst, w4_rsci_adra_d, w4_rsci_ena_d, w4_rsci_qa_d, w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, w4_rsci_oswt, w4_rsci_ena_d_core_psct, w4_rsci_qa_d_mxwt,
      w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct, w4_rsci_adra_d_core_psct_pff,
      w4_rsci_oswt_pff, w4_rsci_adra_d_core_pff
);
  input clk;
  input rst;
  output [23:0] w4_rsci_adra_d;
  output [1:0] w4_rsci_ena_d;
  input [35:0] w4_rsci_qa_d;
  output [1:0] w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input w4_rsci_oswt;
  input [1:0] w4_rsci_ena_d_core_psct;
  output [35:0] w4_rsci_qa_d_mxwt;
  input [1:0] w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input [1:0] w4_rsci_adra_d_core_psct_pff;
  input w4_rsci_oswt_pff;
  input [23:0] w4_rsci_adra_d_core_pff;


  // Interconnect Declarations
  wire w4_rsci_biwt;
  wire w4_rsci_bdwt;
  wire [1:0] w4_rsci_ena_d_core_sct;
  wire [1:0] w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire [23:0] w4_rsci_adra_d_reg;
  wire [1:0] w4_rsci_adra_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [23:0] nl_mnist_mlp_core_w4_rsci_1_w4_rsc_wait_dp_inst_w4_rsci_adra_d_core_pff;
  assign nl_mnist_mlp_core_w4_rsci_1_w4_rsc_wait_dp_inst_w4_rsci_adra_d_core_pff
      = {1'b1 , (w4_rsci_adra_d_core_pff[22:12]) , 1'b0 , (w4_rsci_adra_d_core_pff[10:0])};
  mnist_mlp_core_w4_rsci_1_w4_rsc_wait_ctrl mnist_mlp_core_w4_rsci_1_w4_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .w4_rsci_oswt(w4_rsci_oswt),
      .w4_rsci_ena_d_core_psct(w4_rsci_ena_d_core_psct),
      .w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .w4_rsci_biwt(w4_rsci_biwt),
      .w4_rsci_bdwt(w4_rsci_bdwt),
      .w4_rsci_ena_d_core_sct(w4_rsci_ena_d_core_sct),
      .w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .w4_rsci_adra_d_core_sct_pff(w4_rsci_adra_d_core_sct_iff),
      .w4_rsci_adra_d_core_psct_pff(w4_rsci_adra_d_core_psct_pff),
      .w4_rsci_oswt_pff(w4_rsci_oswt_pff)
    );
  mnist_mlp_core_w4_rsci_1_w4_rsc_wait_dp mnist_mlp_core_w4_rsci_1_w4_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .w4_rsci_adra_d(w4_rsci_adra_d_reg),
      .w4_rsci_qa_d(w4_rsci_qa_d),
      .w4_rsci_qa_d_mxwt(w4_rsci_qa_d_mxwt),
      .w4_rsci_biwt(w4_rsci_biwt),
      .w4_rsci_bdwt(w4_rsci_bdwt),
      .w4_rsci_adra_d_core_sct_pff(w4_rsci_adra_d_core_sct_iff),
      .w4_rsci_adra_d_core_pff(nl_mnist_mlp_core_w4_rsci_1_w4_rsc_wait_dp_inst_w4_rsci_adra_d_core_pff[23:0])
    );
  assign w4_rsci_adra_d = w4_rsci_adra_d_reg;
  assign w4_rsci_ena_d = w4_rsci_ena_d_core_sct;
  assign w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_w2_rsci_1
// ------------------------------------------------------------------


module mnist_mlp_core_w2_rsci_1 (
  clk, rst, w2_rsci_adra_d, w2_rsci_ena_d, w2_rsci_qa_d, w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, w2_rsci_oswt, w2_rsci_adra_d_core_psct, w2_rsci_ena_d_core_psct,
      w2_rsci_qa_d_mxwt, w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct, w2_rsci_adra_d_core_pff,
      w2_rsci_oswt_pff
);
  input clk;
  input rst;
  output [31:0] w2_rsci_adra_d;
  output [1:0] w2_rsci_ena_d;
  input [35:0] w2_rsci_qa_d;
  output [1:0] w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input w2_rsci_oswt;
  input [1:0] w2_rsci_adra_d_core_psct;
  input [1:0] w2_rsci_ena_d_core_psct;
  output [35:0] w2_rsci_qa_d_mxwt;
  input [1:0] w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input [31:0] w2_rsci_adra_d_core_pff;
  input w2_rsci_oswt_pff;


  // Interconnect Declarations
  wire w2_rsci_biwt;
  wire w2_rsci_bdwt;
  wire [1:0] w2_rsci_adra_d_core_sct;
  wire [1:0] w2_rsci_ena_d_core_sct;
  wire [1:0] w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire [31:0] w2_rsci_adra_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_mnist_mlp_core_w2_rsci_1_w2_rsc_wait_dp_inst_w2_rsci_adra_d_core_pff;
  assign nl_mnist_mlp_core_w2_rsci_1_w2_rsc_wait_dp_inst_w2_rsci_adra_d_core_pff
      = {(w2_rsci_adra_d_core_pff[31:16]) , 1'b0 , (w2_rsci_adra_d_core_pff[14:0])};
  mnist_mlp_core_w2_rsci_1_w2_rsc_wait_ctrl mnist_mlp_core_w2_rsci_1_w2_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .w2_rsci_oswt(w2_rsci_oswt),
      .w2_rsci_adra_d_core_psct(w2_rsci_adra_d_core_psct),
      .w2_rsci_ena_d_core_psct(w2_rsci_ena_d_core_psct),
      .w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .w2_rsci_biwt(w2_rsci_biwt),
      .w2_rsci_bdwt(w2_rsci_bdwt),
      .w2_rsci_adra_d_core_sct(w2_rsci_adra_d_core_sct),
      .w2_rsci_ena_d_core_sct(w2_rsci_ena_d_core_sct),
      .w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .w2_rsci_oswt_pff(w2_rsci_oswt_pff)
    );
  mnist_mlp_core_w2_rsci_1_w2_rsc_wait_dp mnist_mlp_core_w2_rsci_1_w2_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .w2_rsci_adra_d(w2_rsci_adra_d_reg),
      .w2_rsci_qa_d(w2_rsci_qa_d),
      .w2_rsci_qa_d_mxwt(w2_rsci_qa_d_mxwt),
      .w2_rsci_biwt(w2_rsci_biwt),
      .w2_rsci_bdwt(w2_rsci_bdwt),
      .w2_rsci_adra_d_core_sct(w2_rsci_adra_d_core_sct),
      .w2_rsci_adra_d_core_pff(nl_mnist_mlp_core_w2_rsci_1_w2_rsc_wait_dp_inst_w2_rsci_adra_d_core_pff[31:0])
    );
  assign w2_rsci_adra_d = w2_rsci_adra_d_reg;
  assign w2_rsci_ena_d = w2_rsci_ena_d_core_sct;
  assign w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_const_size_out_1_rsci
// ------------------------------------------------------------------


module mnist_mlp_core_const_size_out_1_rsci (
  clk, rst, const_size_out_1_rsc_dat, const_size_out_1_rsc_vld, const_size_out_1_rsc_rdy,
      core_wen, const_size_out_1_rsci_oswt, const_size_out_1_rsci_wen_comp
);
  input clk;
  input rst;
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  input const_size_out_1_rsc_rdy;
  input core_wen;
  input const_size_out_1_rsci_oswt;
  output const_size_out_1_rsci_wen_comp;


  // Interconnect Declarations
  wire const_size_out_1_rsci_irdy;
  wire const_size_out_1_rsci_biwt;
  wire const_size_out_1_rsci_bdwt;
  wire const_size_out_1_rsci_bcwt;
  wire const_size_out_1_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd4),
  .width(32'sd16)) const_size_out_1_rsci (
      .irdy(const_size_out_1_rsci_irdy),
      .ivld(const_size_out_1_rsci_ivld_core_sct),
      .idat(16'b0000000000001010),
      .rdy(const_size_out_1_rsc_rdy),
      .vld(const_size_out_1_rsc_vld),
      .dat(const_size_out_1_rsc_dat)
    );
  mnist_mlp_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl mnist_mlp_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .const_size_out_1_rsci_oswt(const_size_out_1_rsci_oswt),
      .const_size_out_1_rsci_irdy(const_size_out_1_rsci_irdy),
      .const_size_out_1_rsci_biwt(const_size_out_1_rsci_biwt),
      .const_size_out_1_rsci_bdwt(const_size_out_1_rsci_bdwt),
      .const_size_out_1_rsci_bcwt(const_size_out_1_rsci_bcwt),
      .const_size_out_1_rsci_ivld_core_sct(const_size_out_1_rsci_ivld_core_sct)
    );
  mnist_mlp_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_dp mnist_mlp_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .const_size_out_1_rsci_oswt(const_size_out_1_rsci_oswt),
      .const_size_out_1_rsci_wen_comp(const_size_out_1_rsci_wen_comp),
      .const_size_out_1_rsci_biwt(const_size_out_1_rsci_biwt),
      .const_size_out_1_rsci_bdwt(const_size_out_1_rsci_bdwt),
      .const_size_out_1_rsci_bcwt(const_size_out_1_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_const_size_in_1_rsci
// ------------------------------------------------------------------


module mnist_mlp_core_const_size_in_1_rsci (
  clk, rst, const_size_in_1_rsc_dat, const_size_in_1_rsc_vld, const_size_in_1_rsc_rdy,
      core_wen, const_size_in_1_rsci_oswt, const_size_in_1_rsci_wen_comp
);
  input clk;
  input rst;
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  input const_size_in_1_rsc_rdy;
  input core_wen;
  input const_size_in_1_rsci_oswt;
  output const_size_in_1_rsci_wen_comp;


  // Interconnect Declarations
  wire const_size_in_1_rsci_irdy;
  wire const_size_in_1_rsci_biwt;
  wire const_size_in_1_rsci_bdwt;
  wire const_size_in_1_rsci_bcwt;
  wire const_size_in_1_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd3),
  .width(32'sd16)) const_size_in_1_rsci (
      .irdy(const_size_in_1_rsci_irdy),
      .ivld(const_size_in_1_rsci_ivld_core_sct),
      .idat(16'b0000001100010000),
      .rdy(const_size_in_1_rsc_rdy),
      .vld(const_size_in_1_rsc_vld),
      .dat(const_size_in_1_rsc_dat)
    );
  mnist_mlp_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl mnist_mlp_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .const_size_in_1_rsci_oswt(const_size_in_1_rsci_oswt),
      .const_size_in_1_rsci_irdy(const_size_in_1_rsci_irdy),
      .const_size_in_1_rsci_biwt(const_size_in_1_rsci_biwt),
      .const_size_in_1_rsci_bdwt(const_size_in_1_rsci_bdwt),
      .const_size_in_1_rsci_bcwt(const_size_in_1_rsci_bcwt),
      .const_size_in_1_rsci_ivld_core_sct(const_size_in_1_rsci_ivld_core_sct)
    );
  mnist_mlp_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_dp mnist_mlp_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .const_size_in_1_rsci_oswt(const_size_in_1_rsci_oswt),
      .const_size_in_1_rsci_wen_comp(const_size_in_1_rsci_wen_comp),
      .const_size_in_1_rsci_biwt(const_size_in_1_rsci_biwt),
      .const_size_in_1_rsci_bdwt(const_size_in_1_rsci_bdwt),
      .const_size_in_1_rsci_bcwt(const_size_in_1_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_layer7_out_rsci
// ------------------------------------------------------------------


module mnist_mlp_core_layer7_out_rsci (
  clk, rst, layer7_out_rsc_dat, layer7_out_rsc_vld, layer7_out_rsc_rdy, core_wen,
      layer7_out_rsci_oswt, layer7_out_rsci_wen_comp, layer7_out_rsci_idat
);
  input clk;
  input rst;
  output [179:0] layer7_out_rsc_dat;
  output layer7_out_rsc_vld;
  input layer7_out_rsc_rdy;
  input core_wen;
  input layer7_out_rsci_oswt;
  output layer7_out_rsci_wen_comp;
  input [179:0] layer7_out_rsci_idat;


  // Interconnect Declarations
  wire layer7_out_rsci_irdy;
  wire layer7_out_rsci_biwt;
  wire layer7_out_rsci_bdwt;
  wire layer7_out_rsci_bcwt;
  wire layer7_out_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  wire [179:0] nl_layer7_out_rsci_idat;
  assign nl_layer7_out_rsci_idat = {6'b000000 , (layer7_out_rsci_idat[173:162]) ,
      6'b000000 , (layer7_out_rsci_idat[155:144]) , 6'b000000 , (layer7_out_rsci_idat[137:126])
      , 6'b000000 , (layer7_out_rsci_idat[119:108]) , 6'b000000 , (layer7_out_rsci_idat[101:90])
      , 6'b000000 , (layer7_out_rsci_idat[83:72]) , 6'b000000 , (layer7_out_rsci_idat[65:54])
      , 6'b000000 , (layer7_out_rsci_idat[47:36]) , 6'b000000 , (layer7_out_rsci_idat[29:18])
      , 6'b000000 , (layer7_out_rsci_idat[11:0])};
  ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd180)) layer7_out_rsci (
      .irdy(layer7_out_rsci_irdy),
      .ivld(layer7_out_rsci_ivld_core_sct),
      .idat(nl_layer7_out_rsci_idat[179:0]),
      .rdy(layer7_out_rsc_rdy),
      .vld(layer7_out_rsc_vld),
      .dat(layer7_out_rsc_dat)
    );
  mnist_mlp_core_layer7_out_rsci_layer7_out_rsc_wait_ctrl mnist_mlp_core_layer7_out_rsci_layer7_out_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .layer7_out_rsci_oswt(layer7_out_rsci_oswt),
      .layer7_out_rsci_irdy(layer7_out_rsci_irdy),
      .layer7_out_rsci_biwt(layer7_out_rsci_biwt),
      .layer7_out_rsci_bdwt(layer7_out_rsci_bdwt),
      .layer7_out_rsci_bcwt(layer7_out_rsci_bcwt),
      .layer7_out_rsci_ivld_core_sct(layer7_out_rsci_ivld_core_sct)
    );
  mnist_mlp_core_layer7_out_rsci_layer7_out_rsc_wait_dp mnist_mlp_core_layer7_out_rsci_layer7_out_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .layer7_out_rsci_oswt(layer7_out_rsci_oswt),
      .layer7_out_rsci_wen_comp(layer7_out_rsci_wen_comp),
      .layer7_out_rsci_biwt(layer7_out_rsci_biwt),
      .layer7_out_rsci_bdwt(layer7_out_rsci_bdwt),
      .layer7_out_rsci_bcwt(layer7_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core_input1_rsci
// ------------------------------------------------------------------


module mnist_mlp_core_input1_rsci (
  clk, rst, input1_rsc_dat, input1_rsc_vld, input1_rsc_rdy, core_wen, input1_rsci_oswt,
      input1_rsci_wen_comp, input1_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [14111:0] input1_rsc_dat;
  input input1_rsc_vld;
  output input1_rsc_rdy;
  input core_wen;
  input input1_rsci_oswt;
  output input1_rsci_wen_comp;
  output [14111:0] input1_rsci_idat_mxwt;


  // Interconnect Declarations
  wire input1_rsci_biwt;
  wire input1_rsci_bdwt;
  wire input1_rsci_bcwt;
  wire input1_rsci_irdy_core_sct;
  wire input1_rsci_ivld;
  wire [14111:0] input1_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd14112)) input1_rsci (
      .rdy(input1_rsc_rdy),
      .vld(input1_rsc_vld),
      .dat(input1_rsc_dat),
      .irdy(input1_rsci_irdy_core_sct),
      .ivld(input1_rsci_ivld),
      .idat(input1_rsci_idat)
    );
  mnist_mlp_core_input1_rsci_input1_rsc_wait_ctrl mnist_mlp_core_input1_rsci_input1_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .input1_rsci_oswt(input1_rsci_oswt),
      .input1_rsci_biwt(input1_rsci_biwt),
      .input1_rsci_bdwt(input1_rsci_bdwt),
      .input1_rsci_bcwt(input1_rsci_bcwt),
      .input1_rsci_irdy_core_sct(input1_rsci_irdy_core_sct),
      .input1_rsci_ivld(input1_rsci_ivld)
    );
  mnist_mlp_core_input1_rsci_input1_rsc_wait_dp mnist_mlp_core_input1_rsci_input1_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input1_rsci_oswt(input1_rsci_oswt),
      .input1_rsci_wen_comp(input1_rsci_wen_comp),
      .input1_rsci_idat_mxwt(input1_rsci_idat_mxwt),
      .input1_rsci_biwt(input1_rsci_biwt),
      .input1_rsci_bdwt(input1_rsci_bdwt),
      .input1_rsci_bcwt(input1_rsci_bcwt),
      .input1_rsci_idat(input1_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp_core
// ------------------------------------------------------------------


module mnist_mlp_core (
  clk, rst, input1_rsc_dat, input1_rsc_vld, input1_rsc_rdy, layer7_out_rsc_dat, layer7_out_rsc_vld,
      layer7_out_rsc_rdy, const_size_in_1_rsc_dat, const_size_in_1_rsc_vld, const_size_in_1_rsc_rdy,
      const_size_out_1_rsc_dat, const_size_out_1_rsc_vld, const_size_out_1_rsc_rdy,
      b2_rsc_dat, b4_rsc_dat, b6_rsc_dat, w2_rsci_adra_d, w2_rsci_ena_d, w2_rsci_qa_d,
      w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, w4_rsci_adra_d, w4_rsci_ena_d,
      w4_rsci_qa_d, w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, w6_rsci_adra_d,
      w6_rsci_ena_d, w6_rsci_qa_d, w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d
);
  input clk;
  input rst;
  input [14111:0] input1_rsc_dat;
  input input1_rsc_vld;
  output input1_rsc_rdy;
  output [179:0] layer7_out_rsc_dat;
  output layer7_out_rsc_vld;
  input layer7_out_rsc_rdy;
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  input const_size_in_1_rsc_rdy;
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  input const_size_out_1_rsc_rdy;
  input [1151:0] b2_rsc_dat;
  input [1151:0] b4_rsc_dat;
  input [179:0] b6_rsc_dat;
  output [31:0] w2_rsci_adra_d;
  output [1:0] w2_rsci_ena_d;
  input [35:0] w2_rsci_qa_d;
  output [1:0] w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [23:0] w4_rsci_adra_d;
  output [1:0] w4_rsci_ena_d;
  input [35:0] w4_rsci_qa_d;
  output [1:0] w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [19:0] w6_rsci_adra_d;
  output [1:0] w6_rsci_ena_d;
  input [35:0] w6_rsci_qa_d;
  output [1:0] w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations
  wire core_wen;
  wire core_wten;
  wire input1_rsci_wen_comp;
  wire [14111:0] input1_rsci_idat_mxwt;
  wire layer7_out_rsci_wen_comp;
  wire const_size_in_1_rsci_wen_comp;
  wire const_size_out_1_rsci_wen_comp;
  wire [35:0] w2_rsci_qa_d_mxwt;
  wire [1151:0] b2_rsci_idat;
  wire [35:0] w4_rsci_qa_d_mxwt;
  wire [1151:0] b4_rsci_idat;
  wire [35:0] w6_rsci_qa_d_mxwt;
  wire [179:0] b6_rsci_idat;
  reg [11:0] layer7_out_rsci_idat_173_162;
  reg [11:0] layer7_out_rsci_idat_155_144;
  reg [11:0] layer7_out_rsci_idat_137_126;
  reg [11:0] layer7_out_rsci_idat_119_108;
  reg [11:0] layer7_out_rsci_idat_101_90;
  reg [11:0] layer7_out_rsci_idat_83_72;
  reg [11:0] layer7_out_rsci_idat_65_54;
  reg [11:0] layer7_out_rsci_idat_47_36;
  reg [11:0] layer7_out_rsci_idat_29_18;
  reg [11:0] layer7_out_rsci_idat_11_0;
  wire [7:0] fsm_output;
  wire nnet_softmax_layer6_t_result_t_softmax_config7_for_1_or_tmp;
  wire [2:0] MultLoop_2_1_acc_3_tmp;
  wire [3:0] nl_MultLoop_2_1_acc_3_tmp;
  wire IndexLoop_IndexLoop_nor_tmp;
  wire [5:0] IndexLoop_mux_1_tmp;
  wire and_dcpl;
  wire or_tmp_1;
  wire or_tmp_2;
  wire mux_tmp_2;
  wire or_tmp_48;
  wire mux_tmp_81;
  wire or_tmp_91;
  wire mux_tmp_183;
  wire mux_tmp_184;
  wire or_tmp_196;
  wire or_tmp_231;
  wire mux_tmp_377;
  wire nand_tmp_14;
  wire mux_tmp_419;
  wire and_dcpl_50;
  wire and_dcpl_51;
  wire and_dcpl_53;
  wire and_dcpl_54;
  wire and_dcpl_55;
  wire and_dcpl_56;
  wire and_dcpl_57;
  wire and_dcpl_58;
  wire and_dcpl_59;
  wire and_dcpl_60;
  wire and_dcpl_62;
  wire and_dcpl_64;
  wire and_dcpl_65;
  wire and_dcpl_66;
  wire and_dcpl_70;
  wire and_dcpl_73;
  wire and_dcpl_75;
  wire and_dcpl_77;
  wire and_dcpl_82;
  wire and_dcpl_84;
  wire and_dcpl_87;
  wire or_dcpl_334;
  wire and_dcpl_92;
  wire and_dcpl_93;
  wire and_dcpl_94;
  wire and_dcpl_95;
  wire and_dcpl_99;
  wire and_dcpl_100;
  wire and_dcpl_101;
  wire and_dcpl_103;
  wire and_dcpl_106;
  wire or_dcpl_337;
  wire or_dcpl_338;
  wire or_dcpl_339;
  wire and_dcpl_109;
  wire or_dcpl_340;
  wire or_dcpl_341;
  wire or_dcpl_342;
  wire or_dcpl_343;
  wire and_dcpl_120;
  wire or_dcpl_344;
  wire or_dcpl_345;
  wire or_dcpl_346;
  wire or_dcpl_347;
  wire and_dcpl_131;
  wire or_dcpl_348;
  wire or_dcpl_349;
  wire and_dcpl_143;
  wire or_dcpl_350;
  wire or_dcpl_351;
  wire and_dcpl_154;
  wire and_dcpl_155;
  wire or_dcpl_362;
  wire or_dcpl_363;
  wire or_dcpl_364;
  wire or_dcpl_365;
  wire or_dcpl_366;
  wire or_dcpl_368;
  wire or_dcpl_369;
  wire or_dcpl_370;
  wire or_dcpl_371;
  wire or_dcpl_372;
  wire or_dcpl_373;
  wire or_dcpl_374;
  wire or_dcpl_375;
  wire or_dcpl_376;
  wire or_dcpl_377;
  wire or_dcpl_378;
  wire or_dcpl_379;
  wire or_dcpl_380;
  wire or_dcpl_381;
  wire or_dcpl_382;
  wire or_dcpl_383;
  wire or_dcpl_384;
  wire or_dcpl_385;
  wire or_dcpl_386;
  wire or_dcpl_387;
  wire or_dcpl_388;
  wire or_dcpl_389;
  wire or_dcpl_390;
  wire or_dcpl_391;
  wire or_dcpl_392;
  wire or_dcpl_393;
  wire or_dcpl_394;
  wire or_dcpl_395;
  wire or_dcpl_396;
  wire or_dcpl_397;
  wire or_dcpl_398;
  wire or_dcpl_399;
  wire or_dcpl_400;
  wire or_dcpl_401;
  wire or_dcpl_402;
  wire or_dcpl_403;
  wire or_dcpl_404;
  wire or_dcpl_405;
  wire or_dcpl_406;
  wire or_dcpl_407;
  wire or_dcpl_408;
  wire or_dcpl_409;
  wire or_dcpl_410;
  wire or_dcpl_411;
  wire or_dcpl_412;
  wire or_dcpl_413;
  wire or_dcpl_414;
  wire or_dcpl_415;
  wire or_dcpl_416;
  wire or_dcpl_417;
  wire or_dcpl_418;
  wire or_dcpl_419;
  wire or_dcpl_420;
  wire or_dcpl_421;
  wire or_dcpl_422;
  wire or_dcpl_423;
  wire or_dcpl_424;
  wire or_dcpl_425;
  wire or_dcpl_426;
  wire or_dcpl_427;
  wire or_dcpl_428;
  wire or_dcpl_429;
  wire or_dcpl_430;
  wire or_dcpl_431;
  wire or_dcpl_432;
  wire or_dcpl_433;
  wire or_dcpl_434;
  wire or_dcpl_435;
  wire or_dcpl_436;
  wire or_dcpl_437;
  wire or_dcpl_438;
  wire or_dcpl_439;
  wire or_dcpl_440;
  wire or_dcpl_441;
  wire or_dcpl_442;
  wire or_dcpl_443;
  wire or_dcpl_444;
  wire or_dcpl_445;
  wire or_dcpl_446;
  wire or_dcpl_447;
  wire or_dcpl_448;
  wire and_dcpl_157;
  wire and_dcpl_158;
  wire and_dcpl_159;
  wire and_dcpl_160;
  wire or_dcpl_455;
  wire or_dcpl_465;
  wire or_dcpl_466;
  wire or_dcpl_467;
  wire or_dcpl_469;
  wire or_dcpl_471;
  wire or_dcpl_472;
  wire or_dcpl_481;
  wire or_dcpl_484;
  wire and_dcpl_169;
  wire and_dcpl_171;
  wire and_dcpl_175;
  wire or_dcpl_490;
  wire and_dcpl_176;
  wire and_dcpl_177;
  wire and_dcpl_178;
  wire and_dcpl_179;
  wire and_dcpl_180;
  wire and_dcpl_181;
  wire and_dcpl_185;
  wire and_dcpl_188;
  wire and_dcpl_189;
  wire or_dcpl_492;
  wire or_dcpl_493;
  wire or_dcpl_494;
  wire or_dcpl_495;
  wire and_dcpl_194;
  wire or_tmp_384;
  wire mux_tmp_488;
  wire and_dcpl_197;
  wire and_dcpl_198;
  wire and_dcpl_199;
  wire and_dcpl_200;
  wire and_dcpl_204;
  wire and_dcpl_205;
  wire and_dcpl_206;
  wire and_dcpl_207;
  wire or_dcpl_498;
  wire or_dcpl_499;
  wire or_dcpl_500;
  wire or_dcpl_501;
  wire and_dcpl_210;
  wire mux_tmp_496;
  wire mux_tmp_497;
  wire mux_tmp_498;
  wire mux_tmp_500;
  wire and_dcpl_211;
  wire and_dcpl_212;
  wire and_dcpl_216;
  wire and_dcpl_217;
  wire and_dcpl_218;
  wire and_dcpl_219;
  wire or_dcpl_502;
  wire or_dcpl_503;
  wire or_dcpl_504;
  wire or_dcpl_505;
  wire and_dcpl_223;
  wire and_dcpl_227;
  wire and_dcpl_228;
  wire and_dcpl_229;
  wire or_dcpl_510;
  wire or_dcpl_511;
  wire or_dcpl_512;
  wire or_dcpl_513;
  wire mux_tmp_513;
  wire mux_tmp_515;
  wire mux_tmp_516;
  wire mux_tmp_517;
  wire mux_tmp_519;
  wire mux_tmp_520;
  wire mux_tmp_521;
  wire and_dcpl_234;
  wire and_dcpl_235;
  wire and_dcpl_238;
  wire and_dcpl_239;
  wire or_dcpl_515;
  wire or_dcpl_516;
  wire or_dcpl_517;
  wire mux_tmp_530;
  wire mux_tmp_532;
  wire and_dcpl_246;
  wire and_dcpl_247;
  wire and_dcpl_250;
  wire and_dcpl_251;
  wire and_dcpl_254;
  wire and_dcpl_255;
  wire or_dcpl_518;
  wire mux_tmp_541;
  wire mux_tmp_543;
  wire and_dcpl_261;
  wire and_dcpl_262;
  wire and_dcpl_263;
  wire and_dcpl_266;
  wire or_dcpl_519;
  wire or_dcpl_520;
  wire mux_tmp_549;
  wire mux_tmp_551;
  wire mux_tmp_552;
  wire mux_tmp_553;
  wire mux_tmp_555;
  wire and_dcpl_274;
  wire and_dcpl_277;
  wire or_dcpl_521;
  wire or_dcpl_522;
  wire and_dcpl_283;
  wire or_dcpl_525;
  wire or_dcpl_526;
  wire and_dcpl_295;
  wire or_dcpl_528;
  wire mux_tmp_570;
  wire or_dcpl_529;
  wire and_dcpl_303;
  wire or_dcpl_531;
  wire and_dcpl_309;
  wire and_dcpl_312;
  wire or_dcpl_533;
  wire or_tmp_449;
  wire mux_tmp_586;
  wire mux_tmp_587;
  wire or_dcpl_534;
  wire mux_tmp_594;
  wire or_dcpl_535;
  wire and_dcpl_324;
  wire and_dcpl_325;
  wire and_dcpl_326;
  wire and_dcpl_329;
  wire or_dcpl_536;
  wire or_dcpl_537;
  wire and_dcpl_334;
  wire mux_tmp_620;
  wire mux_tmp_622;
  wire and_dcpl_338;
  wire and_dcpl_339;
  wire or_dcpl_538;
  wire or_dcpl_539;
  wire or_dcpl_540;
  wire and_dcpl_347;
  wire or_dcpl_541;
  wire mux_tmp_634;
  wire mux_tmp_635;
  wire and_dcpl_353;
  wire and_dcpl_354;
  wire and_dcpl_357;
  wire or_dcpl_543;
  wire or_dcpl_544;
  wire mux_tmp_642;
  wire and_dcpl_365;
  wire or_dcpl_545;
  wire mux_tmp_646;
  wire and_dcpl_369;
  wire or_dcpl_546;
  wire and_dcpl_378;
  wire or_dcpl_547;
  wire mux_tmp_657;
  wire or_dcpl_548;
  wire mux_tmp_670;
  wire mux_tmp_678;
  wire mux_tmp_679;
  wire mux_tmp_680;
  wire mux_tmp_691;
  wire mux_tmp_707;
  wire and_dcpl_410;
  wire and_dcpl_415;
  wire or_dcpl_551;
  wire mux_tmp_713;
  wire mux_tmp_722;
  wire mux_tmp_723;
  wire mux_tmp_724;
  wire and_dcpl_424;
  wire and_dcpl_427;
  wire or_dcpl_552;
  wire and_dcpl_430;
  wire mux_tmp_738;
  wire or_dcpl_554;
  wire mux_tmp_742;
  wire and_dcpl_449;
  wire mux_tmp_771;
  wire mux_tmp_772;
  wire mux_tmp_773;
  wire mux_tmp_774;
  wire or_dcpl_556;
  wire and_dcpl_467;
  wire mux_tmp_787;
  wire mux_tmp_806;
  wire mux_tmp_814;
  wire mux_tmp_819;
  wire mux_tmp_820;
  wire and_dcpl_486;
  wire mux_tmp_829;
  wire mux_tmp_830;
  wire mux_tmp_831;
  wire mux_tmp_837;
  wire mux_tmp_845;
  wire or_dcpl_558;
  wire mux_tmp_860;
  wire mux_tmp_861;
  wire or_dcpl_559;
  wire mux_tmp_870;
  wire and_dcpl_509;
  wire or_dcpl_560;
  wire or_dcpl_561;
  wire and_dcpl_517;
  wire and_dcpl_519;
  wire and_dcpl_520;
  wire mux_tmp_909;
  wire mux_tmp_911;
  wire or_dcpl_571;
  wire or_dcpl_572;
  wire or_dcpl_573;
  wire or_dcpl_574;
  wire or_dcpl_575;
  wire or_dcpl_576;
  wire or_dcpl_577;
  wire or_dcpl_578;
  wire or_dcpl_579;
  wire or_dcpl_580;
  wire or_dcpl_581;
  wire or_dcpl_582;
  wire or_dcpl_583;
  wire or_dcpl_584;
  wire or_dcpl_585;
  wire or_dcpl_586;
  wire or_dcpl_587;
  wire or_dcpl_588;
  wire or_dcpl_589;
  wire or_dcpl_590;
  wire or_dcpl_591;
  wire or_dcpl_592;
  wire or_dcpl_593;
  wire or_dcpl_594;
  wire or_dcpl_595;
  wire or_dcpl_596;
  wire or_dcpl_597;
  wire or_dcpl_598;
  wire or_dcpl_599;
  wire or_dcpl_600;
  wire or_dcpl_601;
  wire or_dcpl_602;
  wire mux_tmp_913;
  wire mux_tmp_914;
  wire mux_tmp_915;
  wire mux_tmp_918;
  wire mux_tmp_925;
  wire mux_tmp_926;
  wire and_dcpl_567;
  wire and_dcpl_570;
  wire mux_tmp_928;
  wire and_dcpl_573;
  wire and_dcpl_576;
  wire mux_tmp_930;
  wire and_dcpl_579;
  wire and_dcpl_584;
  wire and_dcpl_587;
  wire and_dcpl_588;
  wire mux_tmp_933;
  wire and_dcpl_590;
  wire and_dcpl_592;
  wire and_dcpl_623;
  wire and_dcpl_624;
  wire and_dcpl_626;
  wire and_dcpl_658;
  wire and_dcpl_659;
  wire and_dcpl_661;
  wire or_dcpl_607;
  wire or_dcpl_611;
  reg [68:0] SUM_EXP_LOOP_acc_11_itm;
  reg IndexLoop_stage_0;
  reg [3:0] InitAccumLoop_2_iacc_3_0_sva;
  reg [5:0] InitAccumLoop_1_iacc_6_0_sva_5_0;
  reg IndexLoop_stage_0_2;
  reg IndexLoop_asn_3_itm_1;
  reg [4:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1;
  reg [2:0] ReuseLoop_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_outidx_const_assign_1_ReuseLoop_2_asn_tmp_3_2_0_psp_sva_1;
  reg MultLoop_2_and_5_itm_1;
  reg nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_out_index_3_0_sva_1_2;
  reg MultLoop_2_and_14_itm_1;
  reg MultLoop_2_and_15_itm_1;
  reg MultLoop_2_MultLoop_2_nor_2_itm_1;
  reg MultLoop_2_and_6_itm_1;
  reg MultLoop_2_and_7_itm_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_63_sva;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_61_1_sva_2;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_60_1_sva_2;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_6_1_sva_2;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_58_1_sva_2;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_59_1_sva_2;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_0_sva_1;
  wire MultLoop_2_and_m1c;
  wire MultLoop_2_nor_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_123_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_125_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_127_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_129_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_131_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_133_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_135_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_137_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_139_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_141_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_143_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_145_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_147_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_149_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_151_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_153_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_155_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_157_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_159_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_161_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_163_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_165_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_167_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_169_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_171_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_173_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_175_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_177_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_179_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_181_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_183_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_185_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_187_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_189_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_191_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_193_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_195_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_197_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_199_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_201_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_203_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_205_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_207_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_209_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_211_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_213_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_215_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_217_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_219_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_221_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_223_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_225_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_227_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_229_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_231_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_233_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_235_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_237_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_239_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_241_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_243_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_245_m1c;
  wire MultLoop_2_and_28_m1c;
  wire and_514_m1c;
  wire and_509_m1c;
  wire and_505_m1c;
  wire and_503_m1c;
  wire and_501_m1c;
  wire and_497_m1c;
  wire and_493_m1c;
  wire and_491_m1c;
  wire and_486_m1c;
  wire and_484_m1c;
  wire and_480_m1c;
  wire and_476_m1c;
  wire and_474_m1c;
  wire and_472_m1c;
  wire and_470_m1c;
  wire and_459_m1c;
  wire and_457_m1c;
  wire and_443_m1c;
  wire and_441_m1c;
  wire and_436_m1c;
  wire and_434_m1c;
  wire and_427_m1c;
  wire and_424_m1c;
  wire and_420_m1c;
  wire and_415_m1c;
  wire and_410_m1c;
  wire and_408_m1c;
  wire and_404_m1c;
  wire and_397_m1c;
  wire and_395_m1c;
  wire and_391_m1c;
  wire and_389_m1c;
  wire and_383_m1c;
  wire and_378_m1c;
  wire and_372_m1c;
  wire and_365_m1c;
  wire and_357_m1c;
  wire and_350_m1c;
  wire and_342_m1c;
  wire and_337_m1c;
  wire and_329_m1c;
  wire and_321_m1c;
  wire and_317_m1c;
  wire and_556_m1c;
  wire and_312_m1c;
  wire and_554_m1c;
  wire and_306_m1c;
  wire and_300_m1c;
  wire and_295_m1c;
  wire and_288_m1c;
  wire and_283_m1c;
  wire and_277_m1c;
  wire and_269_m1c;
  wire and_266_m1c;
  wire and_258_m1c;
  wire and_250_m1c;
  wire and_244_m1c;
  wire and_238_m1c;
  wire and_226_m1c;
  wire and_215_m1c;
  wire and_550_m1c;
  wire MultLoop_2_and_29_m1c;
  wire MultLoop_2_and_30_m1c;
  wire MultLoop_2_and_31_m1c;
  wire or_1419_tmp;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_371_m1c;
  wire MultLoop_2_and_21_m1c;
  wire and_203_m1c;
  wire MultLoop_2_and_20_m1c;
  wire MultLoop_2_and_25_m1c;
  wire or_1420_tmp;
  wire MultLoop_2_and_24_m1c;
  wire MultLoop_2_and_26_m1c;
  wire MultLoop_2_and_23_m1c;
  reg reg_w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_0_cse;
  reg reg_w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_0_cse;
  reg reg_w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_0_cse;
  reg reg_const_size_out_1_rsci_ivld_core_psct_cse;
  reg reg_layer7_out_rsci_ivld_core_psct_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_and_cse;
  wire nnet_softmax_layer6_t_result_t_softmax_config7_for_1_and_cse;
  wire and_817_cse;
  wire or_888_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_65_cse;
  wire nor_306_cse;
  wire or_864_cse;
  wire mux_661_cse;
  wire or_941_cse;
  wire or_1213_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_62_cse;
  wire or_1405_cse;
  wire nand_52_cse;
  wire [16:0] nnet_relu_layer4_t_layer5_t_relu_config5_for_nnet_relu_layer4_t_layer5_t_relu_config5_for_and_cse;
  wire MultLoop_2_and_cse;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_10_18_6_true_AC_TRN_AC_SAT_18_2_AC_TRN_AC_SAT_exp_arr_and_cse;
  wire operator_67_47_false_AC_TRN_AC_WRAP_and_1_cse;
  wire operator_67_47_false_AC_TRN_AC_WRAP_and_5_cse;
  wire or_10_cse;
  wire or_1298_cse;
  wire or_1398_cse;
  wire nor_298_cse;
  wire and_862_cse;
  wire or_381_cse;
  wire mux_456_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_11_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_10_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_9_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_or_8_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_15_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_14_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_13_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_or_9_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_128_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_96_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_97_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_98_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_99_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_100_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_101_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_102_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_103_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_104_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_105_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_106_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_107_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_108_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_109_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_110_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_111_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_112_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_113_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_114_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_115_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_116_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_117_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_118_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_119_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_120_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_121_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_122_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_123_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_124_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_125_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_129_cse;
  wire mux_33_cse;
  wire or_611_cse;
  wire mux_249_cse;
  wire mux_cse;
  wire nor_310_cse;
  wire mux_509_cse;
  wire mux_389_cse;
  wire mux_421_cse;
  wire mux_425_cse;
  wire [31:0] w2_rsci_adra_d_reg;
  wire [1:0] w2_rsci_ena_d_reg;
  wire [1:0] w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire [23:0] w4_rsci_adra_d_reg;
  wire [1:0] w4_rsci_ena_d_reg;
  wire [1:0] w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire [19:0] w6_rsci_adra_d_reg;
  wire and_73_rmff;
  wire [1:0] w6_rsci_ena_d_reg;
  wire [1:0] w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire MultLoop_2_and_5_itm;
  wire MultLoop_2_and_6_itm;
  wire MultLoop_2_and_7_itm;
  wire [90:0] operator_91_21_false_AC_TRN_AC_WRAP_rshift_itm;
  wire [69:0] operator_71_0_false_AC_TRN_AC_WRAP_lshift_itm;
  wire and_dcpl_730;
  wire and_dcpl_737;
  wire and_dcpl_741;
  wire [6:0] z_out;
  wire and_dcpl_756;
  wire and_dcpl_760;
  wire and_dcpl_764;
  wire and_dcpl_768;
  wire [10:0] z_out_2;
  wire [11:0] nl_z_out_2;
  wire and_dcpl_779;
  wire [5:0] z_out_3;
  wire [6:0] nl_z_out_3;
  wire [3:0] z_out_4;
  wire [4:0] nl_z_out_4;
  wire and_dcpl_926;
  wire and_dcpl_949;
  wire [66:0] z_out_9;
  wire and_dcpl_964;
  wire and_dcpl_967;
  wire [70:0] z_out_10;
  wire [71:0] nl_z_out_10;
  wire and_dcpl_979;
  wire [8:0] z_out_11;
  wire [9:0] nl_z_out_11;
  wire and_dcpl_992;
  wire [19:0] z_out_12;
  wire [20:0] nl_z_out_12;
  wire [21:0] z_out_13;
  wire [22:0] nl_z_out_13;
  wire and_dcpl_1163;
  wire [27:0] z_out_17;
  wire signed [35:0] nl_z_out_17;
  wire and_dcpl_1170;
  wire and_dcpl_1175;
  wire and_dcpl_1180;
  wire and_dcpl_1181;
  wire and_dcpl_1184;
  wire and_dcpl_1185;
  wire and_dcpl_1188;
  wire and_dcpl_1190;
  wire and_dcpl_1192;
  wire and_dcpl_1194;
  wire and_dcpl_1197;
  wire and_dcpl_1199;
  wire and_dcpl_1224;
  wire and_dcpl_1228;
  wire [17:0] z_out_20;
  wire [18:0] nl_z_out_20;
  wire [17:0] z_out_21;
  wire [18:0] nl_z_out_21;
  wire and_dcpl_1278;
  wire and_dcpl_1283;
  wire and_dcpl_1285;
  wire and_dcpl_1287;
  wire and_dcpl_1289;
  wire nor_tmp_215;
  wire and_dcpl_1293;
  wire and_dcpl_1294;
  wire and_dcpl_1297;
  wire and_dcpl_1301;
  wire and_dcpl_1302;
  wire nor_tmp_216;
  wire and_dcpl_1304;
  wire and_dcpl_1306;
  wire and_dcpl_1309;
  wire and_dcpl_1313;
  wire and_dcpl_1314;
  wire nor_tmp_217;
  wire and_dcpl_1316;
  wire and_dcpl_1319;
  wire and_dcpl_1323;
  wire and_dcpl_1325;
  wire and_dcpl_1328;
  wire and_dcpl_1331;
  wire and_dcpl_1334;
  wire and_dcpl_1339;
  wire and_dcpl_1342;
  wire and_dcpl_1344;
  wire and_dcpl_1346;
  wire and_dcpl_1349;
  wire and_dcpl_1350;
  wire and_dcpl_1351;
  wire and_dcpl_1353;
  wire and_dcpl_1354;
  wire not_tmp_680;
  wire and_dcpl_1356;
  wire and_dcpl_1359;
  wire and_dcpl_1362;
  wire and_dcpl_1364;
  wire not_tmp_682;
  wire and_dcpl_1366;
  wire and_dcpl_1367;
  wire and_dcpl_1369;
  wire and_dcpl_1371;
  wire and_dcpl_1374;
  wire and_dcpl_1376;
  wire and_dcpl_1378;
  wire and_dcpl_1380;
  wire and_dcpl_1381;
  wire and_dcpl_1383;
  wire and_dcpl_1385;
  wire and_dcpl_1387;
  wire and_dcpl_1389;
  wire and_dcpl_1391;
  wire and_dcpl_1393;
  wire and_dcpl_1395;
  wire and_dcpl_1396;
  wire and_dcpl_1398;
  wire and_dcpl_1399;
  wire and_dcpl_1401;
  wire and_dcpl_1404;
  wire and_dcpl_1406;
  wire and_dcpl_1408;
  wire and_dcpl_1410;
  wire and_dcpl_1412;
  wire and_dcpl_1413;
  wire and_dcpl_1415;
  wire and_dcpl_1417;
  wire and_dcpl_1419;
  wire and_dcpl_1421;
  wire and_dcpl_1423;
  wire and_dcpl_1425;
  wire and_dcpl_1427;
  wire and_dcpl_1429;
  wire and_dcpl_1430;
  wire and_dcpl_1432;
  wire and_dcpl_1434;
  wire and_dcpl_1436;
  wire and_dcpl_1438;
  wire and_dcpl_1440;
  wire and_dcpl_1442;
  wire and_dcpl_1444;
  wire and_dcpl_1445;
  wire and_dcpl_1448;
  wire and_dcpl_1449;
  wire and_dcpl_1451;
  wire and_dcpl_1474;
  wire and_dcpl_1476;
  wire and_dcpl_1483;
  wire [68:0] z_out_24;
  wire [69:0] nl_z_out_24;
  wire [18:0] z_out_25;
  reg [11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_11_0_lpi_2;
  reg [11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_29_18_lpi_2;
  reg [11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_47_36_lpi_2;
  reg [11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_65_54_lpi_2;
  reg [11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_83_72_lpi_2;
  reg [11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_101_90_lpi_2;
  reg [11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_119_108_lpi_2;
  reg [11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_137_126_lpi_2;
  reg [11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_155_144_lpi_2;
  reg [11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_173_162_lpi_2;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_10_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_9_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_8_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_6_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_58_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_59_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_60_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_61_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_1_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_sva_1;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc0_sva;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc1_sva;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc2_sva;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc3_sva;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc4_sva;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc5_sva;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc6_sva;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc7_sva;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc8_sva;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc9_sva;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc10_sva;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc11_sva;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc12_sva;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc13_sva;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc15_sva;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc14_sva_1;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc13_sva_1;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc12_sva_1;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc11_sva_1;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc10_sva_1;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc9_sva_1;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc8_sva_1;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc7_sva_1;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc6_sva_1;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc5_sva_1;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc4_sva_1;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc3_sva_1;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc2_sva_1;
  reg [5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc1_sva_1;
  reg [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_16_0_lpi_1_dfm;
  reg [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_16_0_lpi_1_dfm;
  reg [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_16_0_lpi_1_dfm;
  reg [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_16_0_lpi_1_dfm;
  reg [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_16_0_lpi_1_dfm;
  reg [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_16_0_lpi_1_dfm;
  reg [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_16_0_lpi_1_dfm;
  reg [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_16_0_lpi_1_dfm;
  reg [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_16_0_lpi_1_dfm;
  reg [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_16_0_lpi_1_dfm;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_31_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_32_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_30_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_33_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_29_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_34_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_28_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_35_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_27_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_36_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_26_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_37_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_25_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_38_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_24_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_39_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_23_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_40_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_22_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_41_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_21_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_42_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_20_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_43_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_19_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_44_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_18_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_45_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_17_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_46_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_16_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_47_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_15_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_48_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_14_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_49_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_13_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_50_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_12_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_51_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_11_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_52_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_10_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_53_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_9_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_54_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_8_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_55_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_7_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_56_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_6_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_57_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_5_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_58_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_4_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_59_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_3_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_60_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_2_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_61_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_62_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_4_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_5_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_3_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_6_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_2_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_7_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_1_sva_1;
  reg [17:0] nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_8_sva_1;
  reg nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_5_sva;
  reg nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_6_sva;
  reg nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_7_sva;
  reg nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_8_sva;
  reg nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_9_sva;
  reg nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_sva;
  reg [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_10_18_6_true_AC_TRN_AC_SAT_18_2_AC_TRN_AC_SAT_exp_arr_0_sva;
  reg [66:0] CALC_EXP_LOOP_2_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva;
  reg [66:0] CALC_EXP_LOOP_3_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva;
  reg [66:0] CALC_EXP_LOOP_4_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva;
  reg [66:0] CALC_EXP_LOOP_5_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva;
  reg [66:0] CALC_EXP_LOOP_6_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva;
  reg [66:0] CALC_EXP_LOOP_7_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva;
  reg [66:0] CALC_EXP_LOOP_8_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva;
  reg [66:0] CALC_EXP_LOOP_9_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva;
  reg [66:0] CALC_EXP_LOOP_10_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva;
  reg [90:0] ac_math_ac_reciprocal_pwl_AC_TRN_71_51_false_AC_TRN_AC_WRAP_91_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1_dfm;
  reg [67:0] SUM_EXP_LOOP_acc_9_itm;
  wire layer7_out_rsci_idat_11_0_mx0c1;
  wire layer7_out_rsci_idat_29_18_mx0c1;
  wire layer7_out_rsci_idat_47_36_mx0c1;
  wire layer7_out_rsci_idat_65_54_mx0c1;
  wire layer7_out_rsci_idat_83_72_mx0c1;
  wire layer7_out_rsci_idat_101_90_mx0c1;
  wire layer7_out_rsci_idat_119_108_mx0c1;
  wire layer7_out_rsci_idat_137_126_mx0c1;
  wire layer7_out_rsci_idat_155_144_mx0c1;
  wire layer7_out_rsci_idat_173_162_mx0c1;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_1_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_61_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_60_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_59_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_58_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_6_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_8_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_9_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_10_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_sva_1_mx2;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_sva_1_mx2;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_sva_2_mx0c3;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_sva_2_mx0c2;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_sva_2_mx0c2;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_sva_2_mx0c2;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_sva_2_mx0c2;
  wire [17:0] InitAccumLoop_2_slc_InitAccumLoop_2_asn_18_17_0_ctmp_sva_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_sva_2_mx0c3;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_sva_2_mx0c3;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_sva_2_mx0c3;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_sva_2_mx0c3;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_sva_2_mx0c3;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_2_mx0c0;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_2_mx0c3;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_2_mx0c4;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_2_mx0c5;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_2_mx0c0;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_2_mx0c4;
  wire [17:0] InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1;
  wire MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_mx0c2;
  wire [17:0] InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1;
  wire [17:0] MultLoop_1_slc_input1_18_17_0_cse_sva_1;
  wire [6:0] IndexLoop_if_acc_4_psp_sva_1;
  wire [7:0] nl_IndexLoop_if_acc_4_psp_sva_1;
  wire [7:0] IndexLoop_if_acc_3_psp_1_sva_1;
  wire [8:0] nl_IndexLoop_if_acc_3_psp_1_sva_1;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_16_0_lpi_1_dfm_mx0w2;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_16_0_lpi_1_dfm_mx0w2;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_16_0_lpi_1_dfm_mx0w2;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_16_0_lpi_1_dfm_mx0w2;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_16_0_lpi_1_dfm_mx0w2;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_16_0_lpi_1_dfm_mx0w2;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire [16:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_16_0_lpi_1_dfm_mx0w0;
  wire nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_4_sva_mx0w1;
  wire nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_3_sva_mx0w1;
  wire nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_2_sva_mx0w1;
  wire nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_sva_mx0w0;
  wire nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_9_sva_mx0w0;
  wire nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_8_sva_mx0w0;
  wire nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_7_sva_mx0w0;
  wire nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_6_sva_mx0w0;
  wire nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_5_sva_mx0w0;
  wire [14:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_1_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_psp_sva_1;
  wire nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_1_sva_1;
  wire [11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000;
  wire [14:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_3_14_0;
  wire [9:0] ROM_1i3_1o10_bb905e8578f158e8f5b59add1dc96bdb2f_1;
  wire [4:0] ROM_1i11_1o5_b94ddd86102738ded3ce1c444a799cda31_1;
  wire [2:0] ROM_1i9_1o3_2fa806bf16b3e0d54016201674d036b62f_1;
  wire [7:0] ROM_1i3_1o8_bdb5a3eca137308489a677a1241b230a2e_1;
  wire [6:0] libraries_leading_sign_71_0_e5d4bd9dc928fda5adf5bf26ec9a2550b9a2_1;
  wire [11:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_conc_231_itm_11_0;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_127_tmp;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_126_tmp;
  wire or_1084_tmp;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_385_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_383_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_381_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_379_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_377_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_375_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_373_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_371_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_369_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_367_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_365_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_363_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_361_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_359_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_357_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_355_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_353_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_351_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_349_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_347_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_345_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_343_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_341_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_339_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_337_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_335_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_333_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_331_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_329_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_327_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_325_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_263_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_57_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_53_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_49_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_45_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_41_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_37_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_33_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_29_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_272_rgt;
  wire MultLoop_and_251_rgt;
  wire MultLoop_and_252_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_243_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_642_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_271_rgt;
  wire MultLoop_and_243_rgt;
  wire MultLoop_and_244_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_637_rgt;
  wire and_225_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_304_rgt;
  wire MultLoop_and_242_rgt;
  wire and_232_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_270_rgt;
  wire MultLoop_and_239_rgt;
  wire MultLoop_and_240_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_630_rgt;
  wire and_243_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_303_rgt;
  wire MultLoop_and_238_rgt;
  wire and_246_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_269_rgt;
  wire MultLoop_and_235_rgt;
  wire MultLoop_and_236_rgt;
  wire and_254_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_268_rgt;
  wire MultLoop_and_233_rgt;
  wire MultLoop_and_234_rgt;
  wire and_261_rgt;
  wire and_265_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_302_rgt;
  wire MultLoop_and_232_rgt;
  wire and_268_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_301_rgt;
  wire MultLoop_and_230_rgt;
  wire and_274_rgt;
  wire and_276_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_300_rgt;
  wire MultLoop_and_228_rgt;
  wire and_280_rgt;
  wire and_282_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_299_rgt;
  wire MultLoop_and_226_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_608_rgt;
  wire and_287_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_298_rgt;
  wire MultLoop_and_224_rgt;
  wire and_292_rgt;
  wire and_294_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_297_rgt;
  wire MultLoop_and_222_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_601_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_267_rgt;
  wire MultLoop_and_219_rgt;
  wire MultLoop_and_220_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_596_rgt;
  wire and_305_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_296_rgt;
  wire MultLoop_and_218_rgt;
  wire and_308_rgt;
  wire and_311_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_295_rgt;
  wire MultLoop_and_214_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_587_rgt;
  wire and_316_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_294_rgt;
  wire MultLoop_and_210_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_582_rgt;
  wire and_320_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_293_rgt;
  wire MultLoop_and_208_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_577_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_266_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_307_rgt;
  wire MultLoop_and_206_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_566_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_571_rgt;
  wire and_334_rgt;
  wire and_336_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_292_rgt;
  wire MultLoop_and_204_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_265_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_306_rgt;
  wire MultLoop_and_202_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_558_rgt;
  wire and_347_rgt;
  wire and_349_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_291_rgt;
  wire MultLoop_and_200_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_552_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_264_rgt;
  wire MultLoop_and_197_rgt;
  wire MultLoop_and_198_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_546_rgt;
  wire and_363_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_263_rgt;
  wire MultLoop_and_195_rgt;
  wire MultLoop_and_196_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_540_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_262_rgt;
  wire MultLoop_and_193_rgt;
  wire MultLoop_and_194_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_534_rgt;
  wire and_376_rgt;
  wire and_377_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_290_rgt;
  wire MultLoop_and_192_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_528_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_261_rgt;
  wire MultLoop_and_189_rgt;
  wire MultLoop_and_190_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_522_rgt;
  wire and_387_rgt;
  wire and_388_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_289_rgt;
  wire MultLoop_and_188_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_260_rgt;
  wire MultLoop_and_185_rgt;
  wire MultLoop_and_186_rgt;
  wire and_393_rgt;
  wire and_394_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_288_rgt;
  wire MultLoop_and_184_rgt;
  wire and_403_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_287_rgt;
  wire MultLoop_and_180_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_258_rgt;
  wire MultLoop_and_177_rgt;
  wire MultLoop_and_178_rgt;
  wire and_409_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_286_rgt;
  wire MultLoop_and_176_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_257_rgt;
  wire MultLoop_and_173_rgt;
  wire MultLoop_and_174_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_480_rgt;
  wire and_419_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_285_rgt;
  wire MultLoop_and_172_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_256_rgt;
  wire MultLoop_and_169_rgt;
  wire MultLoop_and_170_rgt;
  wire and_426_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_284_rgt;
  wire MultLoop_and_168_rgt;
  wire and_430_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_255_rgt;
  wire MultLoop_and_165_rgt;
  wire MultLoop_and_166_rgt;
  wire and_435_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_283_rgt;
  wire MultLoop_and_164_rgt;
  wire and_438_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_254_rgt;
  wire MultLoop_and_161_rgt;
  wire MultLoop_and_162_rgt;
  wire and_442_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_282_rgt;
  wire MultLoop_and_160_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_253_rgt;
  wire MultLoop_and_157_rgt;
  wire MultLoop_and_158_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_252_rgt;
  wire MultLoop_and_155_rgt;
  wire MultLoop_and_156_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_440_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_251_rgt;
  wire MultLoop_and_153_rgt;
  wire MultLoop_and_154_rgt;
  wire and_471_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_281_rgt;
  wire MultLoop_and_152_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_250_rgt;
  wire MultLoop_and_149_rgt;
  wire MultLoop_and_150_rgt;
  wire and_475_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_280_rgt;
  wire MultLoop_and_148_rgt;
  wire and_478_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_249_rgt;
  wire MultLoop_and_145_rgt;
  wire MultLoop_and_146_rgt;
  wire and_482_rgt;
  wire and_483_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_279_rgt;
  wire MultLoop_and_144_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_248_rgt;
  wire MultLoop_and_141_rgt;
  wire MultLoop_and_142_rgt;
  wire and_489_rgt;
  wire and_490_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_278_rgt;
  wire MultLoop_and_140_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_247_rgt;
  wire MultLoop_and_137_rgt;
  wire MultLoop_and_138_rgt;
  wire and_495_rgt;
  wire and_496_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_277_rgt;
  wire MultLoop_and_136_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_397_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_246_rgt;
  wire MultLoop_and_133_rgt;
  wire MultLoop_and_134_rgt;
  wire and_502_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_276_rgt;
  wire MultLoop_and_132_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_245_rgt;
  wire MultLoop_and_129_rgt;
  wire MultLoop_and_130_rgt;
  wire and_507_rgt;
  wire and_508_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_275_rgt;
  wire MultLoop_and_128_rgt;
  wire and_512_rgt;
  wire and_513_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_274_rgt;
  wire MultLoop_and_126_rgt;
  wire and_516_rgt;
  wire and_566_rgt;
  wire and_568_rgt;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd;
  reg [9:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd_2;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_1_ftd;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_1_ftd;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_1_ftd;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd_1;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd_1;
  wire nnet_product_input_t_config2_weight_t_config2_accum_t_1_or_1_ssc;
  wire [67:0] SUM_EXP_LOOP_acc_10_sdt;
  wire [68:0] nl_SUM_EXP_LOOP_acc_10_sdt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_641_cse;
  wire [11:0] CALC_SOFTMAX_LOOP_6_or_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_640_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_629_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_639_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_569_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_521_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_527_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_533_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_545_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_551_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_557_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_570_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_576_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_581_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_586_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_595_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_567_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_600_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_636_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_607_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_539_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_439_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_396_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_479_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_591_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_465_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_456_cse;
  wire nand_152_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_121_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_120_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_119_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_118_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_117_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_116_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_1_ftd_1;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_114_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_1_ftd_1;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_112_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_1_ftd_1;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_110_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_1_ftd_1;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_108_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_107_ssc;
  reg [2:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd;
  reg [10:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_106_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_104_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_1_ftd_1;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_102_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_1_ftd_1;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_100_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_1_ftd_1;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_98_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_1_ftd_1;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_96_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_1_ftd_1;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_94_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_92_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_90_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_88_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_86_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_84_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_82_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_80_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_79_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_78_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_77_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_76_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_75_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_73_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_72_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_70_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_68_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_1_ftd_1;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_64_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_1_ftd_1;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_63_ssc;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_63_1_ftd;
  reg [16:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_63_1_ftd_1;
  reg [2:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_1_ftd;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_447_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_472_m1c;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_482_m1c;
  wire [1:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15;
  wire [1:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15;
  wire [10:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_10_0;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_136_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_444_cse;
  wire and_1161_cse;
  wire [9:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_9_0;
  wire and_1173_cse;
  wire and_1175_cse;
  wire and_1178_cse;
  wire and_1180_cse;
  wire and_1183_cse;
  wire and_1185_cse;
  wire and_1187_cse;
  wire and_1189_cse;
  wire and_1193_cse;
  wire and_1195_cse;
  wire and_1270_cse;
  wire and_1273_cse;
  wire and_1276_cse;
  wire and_1279_cse;
  wire and_1282_cse;
  wire and_1284_cse;
  wire and_1286_cse;
  wire and_1288_cse;
  wire and_1134_cse;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_946_rgt;
  wire nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_948_rgt;
  wire [17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_192_rgt;
  wire [16:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_796_rgt;
  wire or_tmp_922;
  wire not_tmp_1409;
  wire [6:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_745_rgt;
  wire not_tmp_1420;
  wire or_tmp_940;
  wire or_tmp_948;
  wire nand_tmp_52;
  wire or_tmp_957;
  wire nand_tmp_53;
  wire [16:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_747_rgt;
  wire [16:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_748_rgt;
  wire [16:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_749_rgt;
  wire nand_tmp_54;
  wire [16:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_778_rgt;
  wire [16:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_776_rgt;
  wire [16:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_774_rgt;
  wire [16:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_772_rgt;
  wire [16:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_770_rgt;
  wire or_tmp_1095;
  wire [14:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_799_rgt;
  wire or_tmp_1115;
  wire [3:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_766_rgt;
  wire nand_tmp_65;
  wire or_tmp_1128;
  wire nand_tmp_66;
  wire or_tmp_1140;
  wire nand_tmp_67;
  wire mux_tmp_1215;
  wire mux_tmp_1216;
  wire [17:0] MultLoop_mux1h_60_rgt;
  wire [17:0] MultLoop_1_mux1h_65_rgt;
  wire [69:0] SUM_EXP_LOOP_mux_1_rgt;
  reg [1:0] SUM_EXP_LOOP_acc_itm_69_68;
  reg [67:0] SUM_EXP_LOOP_acc_itm_67_0;
  reg [11:0] layer3_out_0_16_0_lpi_1_dfm_11_0;
  reg [1:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_16_15;
  reg [14:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_14_0;
  reg [1:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_16_15;
  reg [14:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_14_0;
  reg [1:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_16_15;
  reg [14:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_14_0;
  reg [1:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_16_15;
  reg [14:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_14_0;
  reg [1:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_16_15;
  reg [14:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_14_0;
  reg [1:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_16_15;
  reg [14:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_14_0;
  wire [1:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15;
  wire [14:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0;
  wire [1:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_16_0_lpi_1_dfm_mx0w2_16_15;
  wire [14:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_16_0_lpi_1_dfm_mx0w2_14_0;
  wire [1:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15;
  wire [14:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0;
  wire [1:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15;
  wire [14:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0;
  wire [1:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15;
  wire [14:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0;
  wire [1:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15;
  wire [14:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0;
  reg [5:0] reg_MultLoop_1_mux_64_itm_1_reg;
  reg [11:0] reg_MultLoop_1_mux_64_itm_1_1_reg;
  reg [5:0] reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_reg;
  reg [11:0] reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_1_reg;
  reg [2:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_2_reg;
  reg reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_4_reg;
  reg [2:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_2_reg;
  reg [11:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg;
  reg [4:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_2_reg;
  reg [11:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_3_reg;
  reg [4:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_2_reg;
  reg [11:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_3_reg;
  reg [4:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_2_reg;
  reg [11:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_3_reg;
  reg [4:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_2_reg;
  reg [1:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_4_reg;
  reg [2:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg;
  reg [2:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_1_reg;
  reg [11:0] reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_2_reg;
  wire nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_3_ssc;
  reg [1:0] reg_nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_16_0_lpi_1_dfm_ftd;
  reg [14:0] reg_nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_16_0_lpi_1_dfm_ftd_1;
  wire [1:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_cse_16_15;
  wire [2:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_cse_14_12;
  wire [11:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_cse_11_0;
  wire [4:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12;
  wire [11:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0;
  wire [4:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12;
  wire [11:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0;
  wire [4:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12;
  wire [11:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0;
  wire [4:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12;
  wire [11:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0;
  wire [4:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12;
  wire [11:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0;
  wire [2:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_12;
  wire [11:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0;
  wire [2:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_12;
  wire nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11;
  wire [4:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12;
  wire [1:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_10;
  wire nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_2_ssc;
  reg [4:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_16_0_lpi_1_dfm_16_12;
  reg [11:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_16_0_lpi_1_dfm_11_0;
  wire nor_942_cse;
  wire nor_943_cse;
  wire nor_944_cse;
  wire mux_989_cse;
  wire nor_936_cse;
  wire nor_937_cse;
  wire mux_990_cse;
  wire nor_923_cse;
  wire and_2658_cse;
  wire nor_662_cse;
  wire and_810_cse_1;
  wire nor_654_cse;
  wire nand_209_cse;
  wire or_1637_cse;
  wire nor_647_cse;
  wire and_2654_cse;
  wire nor_646_cse;
  wire nor_642_cse;
  wire nor_610_cse;
  wire nor_622_cse;
  wire or_865_cse_1;
  wire and_2642_cse;
  wire nor_952_cse;
  wire or_1875_cse;
  wire and_2630_cse;
  wire or_647_cse_1;
  wire nand_191_cse;
  wire nor_560_cse;
  wire nor_959_cse;
  wire mux_1243_cse;
  wire and_2631_cse;
  wire nand_198_cse;
  wire and_2650_cse;
  wire or_1479_cse;
  wire nor_668_cse;
  wire nor_586_cse;
  wire or_1800_cse;
  wire nand_210_cse;
  wire or_1286_cse;
  wire or_1876_cse;
  wire and_558_ssc;
  wire and_2617_ssc;
  reg [1:0] layer3_out_0_16_0_lpi_1_dfm_16_15;
  reg [2:0] layer3_out_0_16_0_lpi_1_dfm_14_12;
  wire mux_1162_cse;
  wire and_2657_cse;
  wire nor_649_cse;
  wire mux_1100_cse;
  wire mux_491_itm;
  wire mux_501_itm;
  wire mux_533_itm;
  wire mux_544_itm;
  wire mux_556_itm;
  wire mux_571_itm;
  wire mux_588_itm;
  wire mux_595_itm;
  wire mux_616_itm;
  wire mux_631_itm;
  wire mux_643_itm;
  wire mux_654_itm;
  wire mux_665_itm;
  wire mux_681_itm;
  wire mux_692_itm;
  wire mux_703_itm;
  wire mux_714_itm;
  wire mux_725_itm;
  wire mux_739_itm;
  wire mux_753_itm;
  wire mux_775_itm;
  wire mux_788_itm;
  wire mux_802_itm;
  wire mux_815_itm;
  wire mux_832_itm;
  wire mux_846_itm;
  wire mux_850_itm;
  wire mux_856_itm;
  wire mux_862_itm;
  wire mux_867_itm;
  wire mux_872_itm;
  wire SUM_EXP_LOOP_nor_itm;
  wire ReuseLoop_nor_itm;
  wire ReuseLoop_or_itm;
  wire IndexLoop_if_nor_itm;
  wire operator_18_8_true_AC_TRN_AC_WRAP_1_or_itm;
  wire SUM_EXP_LOOP_nor_2_itm;
  wire ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_10_cse;
  wire nnet_softmax_layer6_t_result_t_softmax_config7_for_3_and_seb;
  wire nnet_softmax_layer6_t_result_t_softmax_config7_for_6_and_seb;
  wire nnet_softmax_layer6_t_result_t_softmax_config7_for_4_and_seb;
  wire nnet_softmax_layer6_t_result_t_softmax_config7_for_5_and_seb;
  wire nnet_softmax_layer6_t_result_t_softmax_config7_for_7_and_seb;
  wire ReuseLoop_and_2_cse;
  wire ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_7_cse;
  wire ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_2_cse;
  wire z_out_1_3;
  wire [147:0] z_out_18_157_10;
  wire [17:0] z_out_19_27_10;
  wire [14:0] z_out_23_22_8;
  wire [14:0] ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_19_cse;
  wire [18:0] ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_sdt;
  wire [19:0] nl_ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_sdt;
  wire and_2670_cse;

  wire[0:0] mux_471_nl;
  wire[0:0] mux_470_nl;
  wire[0:0] or_1411_nl;
  wire[0:0] nand_61_nl;
  wire[0:0] or_713_nl;
  wire[0:0] nor_941_nl;
  wire[5:0] InitAccumLoop_1_iacc_mux_nl;
  wire[0:0] nand_149_nl;
  wire[0:0] mux_478_nl;
  wire[0:0] mux_477_nl;
  wire[0:0] nand_99_nl;
  wire[0:0] mux_152_nl;
  wire[0:0] mux_151_nl;
  wire[0:0] or_378_nl;
  wire[0:0] or_377_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_6_or_1_nl;
  wire[2:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_3_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl;
  wire[2:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_3_nor_2_nl;
  wire[11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_3_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_1_nl;
  wire[11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_3_nor_3_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_644_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_273_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_305_nl;
  wire[0:0] mux_486_nl;
  wire[0:0] or_880_nl;
  wire[0:0] and_193_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_652_nl;
  wire[0:0] and_174_nl;
  wire[0:0] mux_1057_nl;
  wire[0:0] nor_663_nl;
  wire[0:0] mux_1056_nl;
  wire[0:0] mux_1055_nl;
  wire[0:0] mux_1054_nl;
  wire[0:0] or_1553_nl;
  wire[0:0] nand_158_nl;
  wire[0:0] nand_213_nl;
  wire[0:0] or_1548_nl;
  wire[0:0] mux_1053_nl;
  wire[0:0] or_1547_nl;
  wire[0:0] nand_157_nl;
  wire[0:0] mux_1052_nl;
  wire[0:0] nor_666_nl;
  wire[0:0] nor_667_nl;
  wire[0:0] mux_1051_nl;
  wire[0:0] mux_1064_nl;
  wire[0:0] mux_1063_nl;
  wire[0:0] mux_1062_nl;
  wire[0:0] mux_1061_nl;
  wire[0:0] nor_669_nl;
  wire[0:0] and_2660_nl;
  wire[0:0] nor_671_nl;
  wire[0:0] nor_672_nl;
  wire[0:0] mux_1060_nl;
  wire[0:0] or_1561_nl;
  wire[0:0] nand_160_nl;
  wire[0:0] nor_674_nl;
  wire[0:0] mux_1059_nl;
  wire[0:0] mux_1058_nl;
  wire[0:0] nand_159_nl;
  wire[0:0] mux_1071_nl;
  wire[0:0] mux_1070_nl;
  wire[0:0] mux_1069_nl;
  wire[0:0] nor_675_nl;
  wire[0:0] and_2663_nl;
  wire[0:0] mux_1068_nl;
  wire[0:0] mux_1067_nl;
  wire[0:0] nor_676_nl;
  wire[0:0] nor_677_nl;
  wire[0:0] nor_678_nl;
  wire[0:0] mux_1066_nl;
  wire[0:0] mux_1065_nl;
  wire[0:0] nor_679_nl;
  wire[0:0] nor_680_nl;
  wire[0:0] and_2665_nl;
  wire[0:0] nor_682_nl;
  wire[0:0] and_591_nl;
  wire[0:0] and_593_nl;
  wire[0:0] mux_934_nl;
  wire[0:0] and_587_nl;
  wire[0:0] and_588_nl;
  wire[0:0] mux_523_nl;
  wire[0:0] mux_522_nl;
  wire[2:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_6_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl;
  wire[2:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_6_nor_2_nl;
  wire[11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_6_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_1_nl;
  wire[11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_6_nor_3_nl;
  wire[0:0] and_615_nl;
  wire[0:0] and_616_nl;
  wire[0:0] mux_1074_nl;
  wire[0:0] mux_1073_nl;
  wire[0:0] mux_1072_nl;
  wire[0:0] nor_659_nl;
  wire[0:0] nor_660_nl;
  wire[0:0] nor_661_nl;
  wire[0:0] mux_1077_nl;
  wire[0:0] mux_1076_nl;
  wire[0:0] mux_1075_nl;
  wire[0:0] nor_655_nl;
  wire[0:0] nor_656_nl;
  wire[0:0] nor_657_nl;
  wire[0:0] and_638_nl;
  wire[0:0] and_639_nl;
  wire[0:0] and_662_nl;
  wire[0:0] and_664_nl;
  wire[0:0] mux_950_nl;
  wire[0:0] and_685_nl;
  wire[0:0] and_686_nl;
  wire[0:0] and_705_nl;
  wire[0:0] and_709_nl;
  wire[0:0] and_702_nl;
  wire[0:0] and_704_nl;
  wire[0:0] mux_959_nl;
  wire[0:0] and_595_nl;
  wire[0:0] and_596_nl;
  wire[0:0] and_699_nl;
  wire[0:0] and_701_nl;
  wire[0:0] and_696_nl;
  wire[0:0] and_698_nl;
  wire[0:0] mux_958_nl;
  wire[0:0] mux_417_nl;
  wire[0:0] and_693_nl;
  wire[0:0] and_695_nl;
  wire[0:0] and_691_nl;
  wire[0:0] and_692_nl;
  wire[0:0] mux_957_nl;
  wire[0:0] mux_607_nl;
  wire[0:0] mux_606_nl;
  wire[0:0] mux_605_nl;
  wire[0:0] mux_604_nl;
  wire[0:0] mux_603_nl;
  wire[0:0] mux_171_nl;
  wire[0:0] or_870_nl;
  wire[0:0] or_1001_nl;
  wire[0:0] or_649_nl;
  wire[0:0] mux_1082_nl;
  wire[0:0] mux_1081_nl;
  wire[0:0] nand_164_nl;
  wire[0:0] mux_1080_nl;
  wire[0:0] or_1598_nl;
  wire[0:0] or_1596_nl;
  wire[0:0] mux_1079_nl;
  wire[0:0] or_1595_nl;
  wire[0:0] mux_1078_nl;
  wire[0:0] or_1593_nl;
  wire[0:0] mux_1087_nl;
  wire[0:0] mux_1086_nl;
  wire[0:0] and_2656_nl;
  wire[0:0] mux_1085_nl;
  wire[0:0] mux_1084_nl;
  wire[0:0] nor_650_nl;
  wire[0:0] nor_651_nl;
  wire[0:0] mux_1083_nl;
  wire[0:0] nor_652_nl;
  wire[0:0] nor_653_nl;
  wire[9:0] ReuseLoop_ReuseLoop_and_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_470_nl;
  wire[0:0] mux_1091_nl;
  wire[0:0] mux_1090_nl;
  wire[0:0] nor_945_nl;
  wire[0:0] mux_1089_nl;
  wire[0:0] mux_1088_nl;
  wire[0:0] nor_946_nl;
  wire[0:0] nor_947_nl;
  wire[0:0] nor_948_nl;
  wire[0:0] and_689_nl;
  wire[0:0] and_690_nl;
  wire[0:0] mux_623_nl;
  wire[0:0] mux_621_nl;
  wire[0:0] mux_435_nl;
  wire[0:0] and_599_nl;
  wire[0:0] and_600_nl;
  wire[0:0] mux_1099_nl;
  wire[0:0] mux_1098_nl;
  wire[0:0] mux_1097_nl;
  wire[0:0] or_1623_nl;
  wire[0:0] mux_1096_nl;
  wire[0:0] or_1616_nl;
  wire[0:0] mux_1092_nl;
  wire[0:0] mux_1106_nl;
  wire[0:0] mux_1105_nl;
  wire[0:0] mux_1104_nl;
  wire[0:0] or_1632_nl;
  wire[0:0] mux_1103_nl;
  wire[0:0] or_1625_nl;
  wire[0:0] and_687_nl;
  wire[0:0] and_688_nl;
  wire[0:0] mux_956_nl;
  wire[0:0] mux_636_nl;
  wire[0:0] and_601_nl;
  wire[0:0] and_602_nl;
  wire[0:0] mux_1112_nl;
  wire[0:0] mux_1111_nl;
  wire[0:0] and_2651_nl;
  wire[0:0] mux_1110_nl;
  wire[0:0] nor_641_nl;
  wire[0:0] mux_1109_nl;
  wire[0:0] nor_643_nl;
  wire[0:0] nor_644_nl;
  wire[0:0] mux_1108_nl;
  wire[0:0] mux_1107_nl;
  wire[0:0] or_1636_nl;
  wire[0:0] or_1634_nl;
  wire[0:0] mux_1118_nl;
  wire[0:0] mux_1117_nl;
  wire[0:0] nor_645_nl;
  wire[0:0] mux_1116_nl;
  wire[0:0] or_1656_nl;
  wire[0:0] mux_1115_nl;
  wire[0:0] mux_1114_nl;
  wire[0:0] nand_214_nl;
  wire[0:0] or_1652_nl;
  wire[0:0] or_1651_nl;
  wire[0:0] mux_1113_nl;
  wire[0:0] nor_648_nl;
  wire[0:0] and_683_nl;
  wire[0:0] and_684_nl;
  wire[0:0] mux_955_nl;
  wire[0:0] mux_647_nl;
  wire[0:0] and_603_nl;
  wire[0:0] and_604_nl;
  wire[0:0] mux_1124_nl;
  wire[0:0] mux_1123_nl;
  wire[0:0] and_2648_nl;
  wire[0:0] mux_1122_nl;
  wire[0:0] nor_633_nl;
  wire[0:0] and_2649_nl;
  wire[0:0] mux_1121_nl;
  wire[0:0] nor_634_nl;
  wire[0:0] nor_635_nl;
  wire[0:0] nor_636_nl;
  wire[0:0] mux_1120_nl;
  wire[0:0] mux_1119_nl;
  wire[0:0] or_1660_nl;
  wire[0:0] nand_204_nl;
  wire[0:0] mux_1129_nl;
  wire[0:0] mux_1128_nl;
  wire[0:0] nor_637_nl;
  wire[0:0] mux_1127_nl;
  wire[0:0] mux_1126_nl;
  wire[0:0] nor_638_nl;
  wire[0:0] nor_639_nl;
  wire[0:0] nor_640_nl;
  wire[0:0] mux_1125_nl;
  wire[0:0] or_1672_nl;
  wire[0:0] or_1671_nl;
  wire[0:0] and_681_nl;
  wire[0:0] and_682_nl;
  wire[0:0] mux_658_nl;
  wire[0:0] and_605_nl;
  wire[0:0] and_606_nl;
  wire[0:0] mux_1133_nl;
  wire[0:0] nor_954_nl;
  wire[0:0] mux_1132_nl;
  wire[0:0] mux_1131_nl;
  wire[0:0] mux_1130_nl;
  wire[0:0] nor_955_nl;
  wire[0:0] nor_956_nl;
  wire[0:0] nor_957_nl;
  wire[0:0] and_679_nl;
  wire[0:0] and_680_nl;
  wire[0:0] mux_954_nl;
  wire[0:0] mux_671_nl;
  wire[0:0] and_607_nl;
  wire[0:0] and_608_nl;
  wire[0:0] mux_1139_nl;
  wire[0:0] mux_1138_nl;
  wire[0:0] or_1694_nl;
  wire[0:0] mux_1137_nl;
  wire[0:0] or_1688_nl;
  wire[0:0] and_677_nl;
  wire[0:0] and_678_nl;
  wire[0:0] mux_690_nl;
  wire[0:0] or_1083_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_259_nl;
  wire[0:0] MultLoop_and_181_nl;
  wire[0:0] MultLoop_and_182_nl;
  wire[0:0] and_400_nl;
  wire[0:0] and_675_nl;
  wire[0:0] and_676_nl;
  wire[0:0] mux_953_nl;
  wire[0:0] mux_698_nl;
  wire[2:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_4_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl;
  wire[2:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_4_nor_2_nl;
  wire[1:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_4_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_1_nl;
  wire[1:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_4_nor_3_nl;
  wire[9:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_4_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_2_nl;
  wire[9:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_4_nor_4_nl;
  wire[0:0] and_611_nl;
  wire[0:0] and_612_nl;
  wire[0:0] mux_1144_nl;
  wire[0:0] nor_623_nl;
  wire[0:0] mux_1143_nl;
  wire[0:0] mux_1142_nl;
  wire[0:0] and_2647_nl;
  wire[0:0] mux_1141_nl;
  wire[0:0] nor_624_nl;
  wire[0:0] nor_625_nl;
  wire[0:0] mux_1140_nl;
  wire[0:0] nor_626_nl;
  wire[0:0] nor_627_nl;
  wire[0:0] nor_628_nl;
  wire[0:0] mux_1147_nl;
  wire[0:0] and_2644_nl;
  wire[0:0] mux_1146_nl;
  wire[0:0] and_2645_nl;
  wire[0:0] mux_1145_nl;
  wire[0:0] nor_619_nl;
  wire[0:0] nor_620_nl;
  wire[0:0] nor_621_nl;
  wire[0:0] and_673_nl;
  wire[0:0] and_674_nl;
  wire[0:0] mux_708_nl;
  wire[2:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_5_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl;
  wire[2:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_5_nor_2_nl;
  wire[11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_5_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_1_nl;
  wire[11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_5_nor_3_nl;
  wire[0:0] and_613_nl;
  wire[0:0] and_614_nl;
  wire[0:0] mux_1150_nl;
  wire[0:0] mux_1149_nl;
  wire[0:0] nor_615_nl;
  wire[0:0] mux_1148_nl;
  wire[0:0] nor_617_nl;
  wire[0:0] nor_618_nl;
  wire[0:0] mux_1153_nl;
  wire[0:0] mux_1152_nl;
  wire[0:0] mux_1151_nl;
  wire[0:0] nor_611_nl;
  wire[0:0] nor_613_nl;
  wire[0:0] nor_614_nl;
  wire[0:0] and_671_nl;
  wire[0:0] and_672_nl;
  wire[0:0] mux_952_nl;
  wire[0:0] mux_717_nl;
  wire[2:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_7_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl;
  wire[2:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_7_nor_2_nl;
  wire[11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_7_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_1_nl;
  wire[11:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_7_nor_3_nl;
  wire[0:0] and_617_nl;
  wire[0:0] and_618_nl;
  wire[0:0] mux_1157_nl;
  wire[0:0] mux_1156_nl;
  wire[0:0] mux_1155_nl;
  wire[0:0] and_2643_nl;
  wire[0:0] nor_608_nl;
  wire[0:0] mux_1154_nl;
  wire[0:0] nor_609_nl;
  wire[0:0] mux_1160_nl;
  wire[0:0] mux_1159_nl;
  wire[0:0] nor_604_nl;
  wire[0:0] mux_1158_nl;
  wire[0:0] or_1729_nl;
  wire[0:0] or_1728_nl;
  wire[0:0] nor_605_nl;
  wire[0:0] and_669_nl;
  wire[0:0] and_670_nl;
  wire[0:0] mux_729_nl;
  wire[14:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_8_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl;
  wire[14:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_8_nor_2_nl;
  wire[0:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_8_and_nl;
  wire[0:0] and_619_nl;
  wire[0:0] and_620_nl;
  wire[0:0] and_2640_nl;
  wire[0:0] mux_1161_nl;
  wire[0:0] nor_601_nl;
  wire[0:0] nor_602_nl;
  wire[0:0] and_2641_nl;
  wire[0:0] mux_1163_nl;
  wire[0:0] nor_603_nl;
  wire[0:0] mux_1166_nl;
  wire[0:0] and_667_nl;
  wire[0:0] and_668_nl;
  wire[0:0] mux_951_nl;
  wire[0:0] mux_745_nl;
  wire[0:0] mux_744_nl;
  wire[0:0] mux_743_nl;
  wire[14:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_9_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl;
  wire[14:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_9_nor_2_nl;
  wire[0:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_9_and_nl;
  wire[0:0] and_621_nl;
  wire[0:0] and_622_nl;
  wire[0:0] mux_1169_nl;
  wire[0:0] mux_1168_nl;
  wire[0:0] and_2637_nl;
  wire[0:0] mux_1167_nl;
  wire[0:0] nor_594_nl;
  wire[0:0] nor_595_nl;
  wire[0:0] nor_596_nl;
  wire[0:0] nor_597_nl;
  wire[0:0] mux_1173_nl;
  wire[0:0] mux_1172_nl;
  wire[0:0] nor_589_nl;
  wire[0:0] nor_590_nl;
  wire[0:0] mux_1171_nl;
  wire[0:0] mux_1170_nl;
  wire[0:0] nor_591_nl;
  wire[0:0] nor_592_nl;
  wire[0:0] nor_593_nl;
  wire[0:0] and_665_nl;
  wire[0:0] and_666_nl;
  wire[0:0] or_9_nl;
  wire[1:0] MultLoop_1_1_MultLoop_1_mux_nl;
  wire[14:0] IndexLoop_ir_asn_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_3_14_IndexLoop_ir_and_nl;
  wire[14:0] IndexLoop_ir_IndexLoop_ir_mux_nl;
  wire[14:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_10_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl;
  wire[14:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_10_nor_2_nl;
  wire[0:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_10_and_nl;
  wire[0:0] nor_372_nl;
  wire[0:0] mux_887_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] mux_885_nl;
  wire[14:0] MultLoop_1_1_MultLoop_1_mux_1_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_484_nl;
  wire[0:0] mux_1181_nl;
  wire[0:0] mux_1180_nl;
  wire[0:0] mux_1179_nl;
  wire[0:0] or_1771_nl;
  wire[0:0] or_1770_nl;
  wire[0:0] mux_1178_nl;
  wire[0:0] or_1767_nl;
  wire[0:0] mux_1177_nl;
  wire[0:0] mux_1176_nl;
  wire[0:0] mux_1175_nl;
  wire[0:0] or_1763_nl;
  wire[0:0] mux_1174_nl;
  wire[0:0] or_1758_nl;
  wire[0:0] or_1756_nl;
  wire[0:0] mux_1186_nl;
  wire[0:0] mux_1185_nl;
  wire[0:0] mux_1184_nl;
  wire[0:0] mux_1183_nl;
  wire[0:0] nor_583_nl;
  wire[0:0] and_2635_nl;
  wire[0:0] and_2636_nl;
  wire[0:0] mux_1182_nl;
  wire[0:0] nor_585_nl;
  wire[0:0] nor_587_nl;
  wire[0:0] nor_588_nl;
  wire[0:0] and_658_nl;
  wire[0:0] and_659_nl;
  wire[0:0] mux_1191_nl;
  wire[0:0] mux_1190_nl;
  wire[0:0] mux_1189_nl;
  wire[0:0] or_1788_nl;
  wire[0:0] mux_1188_nl;
  wire[0:0] nand_177_nl;
  wire[0:0] mux_1187_nl;
  wire[0:0] or_1786_nl;
  wire[0:0] or_1784_nl;
  wire[0:0] or_1783_nl;
  wire[0:0] mux_1194_nl;
  wire[0:0] nor_578_nl;
  wire[0:0] mux_1193_nl;
  wire[0:0] mux_1192_nl;
  wire[0:0] or_1792_nl;
  wire[0:0] nand_178_nl;
  wire[0:0] nor_580_nl;
  wire[10:0] ReuseLoop_1_ir_ReuseLoop_1_ir_and_nl;
  wire[8:0] ReuseLoop_2_ir_ReuseLoop_2_ir_and_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_446_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_845_nl;
  wire[0:0] and_656_nl;
  wire[0:0] and_657_nl;
  wire[0:0] mux_949_nl;
  wire[0:0] mux_796_nl;
  wire[0:0] and_627_nl;
  wire[0:0] and_629_nl;
  wire[0:0] mux_1198_nl;
  wire[0:0] mux_1197_nl;
  wire[0:0] or_1797_nl;
  wire[0:0] mux_1196_nl;
  wire[0:0] or_1794_nl;
  wire[0:0] and_654_nl;
  wire[0:0] and_655_nl;
  wire[0:0] mux_807_nl;
  wire[0:0] and_630_nl;
  wire[0:0] and_631_nl;
  wire[0:0] mux_1207_nl;
  wire[0:0] mux_1206_nl;
  wire[0:0] or_1803_nl;
  wire[0:0] mux_1205_nl;
  wire[0:0] mux_1204_nl;
  wire[0:0] mux_1203_nl;
  wire[0:0] or_1802_nl;
  wire[0:0] mux_1202_nl;
  wire[0:0] or_1801_nl;
  wire[0:0] mux_1201_nl;
  wire[0:0] mux_1200_nl;
  wire[0:0] mux_1199_nl;
  wire[0:0] or_1799_nl;
  wire[0:0] and_652_nl;
  wire[0:0] and_653_nl;
  wire[0:0] mux_948_nl;
  wire[0:0] mux_822_nl;
  wire[0:0] mux_821_nl;
  wire[0:0] and_632_nl;
  wire[0:0] and_633_nl;
  wire[0:0] mux_1212_nl;
  wire[0:0] mux_1211_nl;
  wire[0:0] or_1809_nl;
  wire[0:0] mux_1210_nl;
  wire[0:0] or_1808_nl;
  wire[0:0] and_650_nl;
  wire[0:0] and_651_nl;
  wire[0:0] mux_838_nl;
  wire[0:0] and_634_nl;
  wire[0:0] and_635_nl;
  wire[0:0] mux_1217_nl;
  wire[0:0] mux_1216_nl;
  wire[0:0] mux_1215_nl;
  wire[0:0] and_648_nl;
  wire[0:0] and_649_nl;
  wire[0:0] mux_947_nl;
  wire[0:0] and_636_nl;
  wire[0:0] and_637_nl;
  wire[0:0] mux_944_nl;
  wire[0:0] and_646_nl;
  wire[0:0] and_647_nl;
  wire[0:0] and_640_nl;
  wire[0:0] and_641_nl;
  wire[0:0] mux_945_nl;
  wire[0:0] and_644_nl;
  wire[0:0] and_645_nl;
  wire[0:0] mux_946_nl;
  wire[0:0] and_642_nl;
  wire[0:0] and_643_nl;
  wire[0:0] IndexLoop_mux1h_9_nl;
  wire[0:0] nnet_dense_large_input_t_layer2_t_config2_if_nnet_dense_large_input_t_layer2_t_config2_if_and_nl;
  wire[0:0] nnet_dense_large_input_t_layer2_t_config2_if_nnet_dense_large_input_t_layer2_t_config2_if_and_1_nl;
  wire[0:0] and_830_nl;
  wire[0:0] IndexLoop_or_1_nl;
  wire[0:0] mux_883_nl;
  wire[0:0] mux_882_nl;
  wire[0:0] or_1413_nl;
  wire[0:0] mux_881_nl;
  wire[0:0] or_1414_nl;
  wire[0:0] or_461_nl;
  wire[0:0] or_1416_nl;
  wire[0:0] mux_688_nl;
  wire[0:0] mux_687_nl;
  wire[5:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_mux_nl;
  wire[5:0] IndexLoop_if_acc_nl;
  wire[6:0] nl_IndexLoop_if_acc_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_and_14_nl;
  wire[0:0] nand_148_nl;
  wire[0:0] mux_890_nl;
  wire[0:0] nor_217_nl;
  wire[0:0] nor_353_nl;
  wire[0:0] mux_10_nl;
  wire[17:0] MultLoop_mux_129_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_63_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_63_nl;
  wire[0:0] MultLoop_and_253_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_185_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_62_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_62_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_372_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_184_nl;
  wire[17:0] MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_30_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_29_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_28_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_27_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_26_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_25_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_24_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_23_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_22_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_21_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_20_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_19_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_18_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_17_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_16_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_15_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_14_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_13_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_12_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_11_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_10_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_9_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_8_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_7_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_6_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_5_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_4_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_3_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_2_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_1_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_63_nl;
  wire[0:0] MultLoop_or_7_nl;
  wire[0:0] MultLoop_or_8_nl;
  wire[0:0] MultLoop_and_250_nl;
  wire[0:0] and_541_nl;
  wire[0:0] MultLoop_and_261_nl;
  wire[0:0] MultLoop_2_and_32_nl;
  wire[0:0] MultLoop_and_262_nl;
  wire[0:0] MultLoop_2_and_37_nl;
  wire[0:0] MultLoop_2_and_39_nl;
  wire[0:0] and_542_nl;
  wire[0:0] mux_892_nl;
  wire[0:0] mux_891_nl;
  wire[0:0] mux_1223_nl;
  wire[0:0] mux_1222_nl;
  wire[0:0] nand_183_nl;
  wire[0:0] mux_1221_nl;
  wire[0:0] or_1820_nl;
  wire[0:0] nand_182_nl;
  wire[0:0] mux_1218_nl;
  wire[0:0] nor_569_nl;
  wire[0:0] nor_570_nl;
  wire[0:0] mux_1227_nl;
  wire[0:0] nor_571_nl;
  wire[0:0] mux_1226_nl;
  wire[0:0] mux_1225_nl;
  wire[0:0] nor_572_nl;
  wire[0:0] nor_573_nl;
  wire[0:0] mux_1224_nl;
  wire[0:0] or_1825_nl;
  wire[17:0] MultLoop_1_mux_64_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_62_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_31_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_32_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_33_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_34_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_35_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_36_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_37_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_38_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_39_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_40_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_41_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_42_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_43_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_44_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_45_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_46_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_47_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_48_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_49_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_50_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_51_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_52_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_53_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_54_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_55_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_56_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_57_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_58_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_59_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_60_nl;
  wire[17:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_61_nl;
  wire[0:0] MultLoop_1_or_3_nl;
  wire[0:0] MultLoop_1_or_4_nl;
  wire[0:0] MultLoop_and_247_nl;
  wire[0:0] and_547_nl;
  wire[0:0] MultLoop_2_and_42_nl;
  wire[0:0] MultLoop_1_and_66_nl;
  wire[0:0] MultLoop_2_and_51_nl;
  wire[0:0] MultLoop_2_and_47_nl;
  wire[0:0] MultLoop_2_and_45_nl;
  wire[0:0] and_552_nl;
  wire[0:0] and_548_nl;
  wire[0:0] mux_901_nl;
  wire[0:0] mux_460_nl;
  wire[0:0] mux_1235_nl;
  wire[0:0] mux_1234_nl;
  wire[0:0] and_2625_nl;
  wire[0:0] nor_558_nl;
  wire[0:0] nor_559_nl;
  wire[0:0] mux_1233_nl;
  wire[0:0] mux_1232_nl;
  wire[0:0] or_1837_nl;
  wire[0:0] mux_1231_nl;
  wire[0:0] nand_192_nl;
  wire[0:0] mux_1230_nl;
  wire[0:0] or_1834_nl;
  wire[0:0] or_1833_nl;
  wire[0:0] nand_185_nl;
  wire[0:0] mux_1229_nl;
  wire[0:0] mux_1228_nl;
  wire[0:0] mux_1241_nl;
  wire[0:0] and_2627_nl;
  wire[0:0] mux_1240_nl;
  wire[0:0] mux_1239_nl;
  wire[0:0] nor_561_nl;
  wire[0:0] and_2628_nl;
  wire[0:0] mux_1238_nl;
  wire[0:0] nor_562_nl;
  wire[0:0] mux_1237_nl;
  wire[0:0] nor_563_nl;
  wire[0:0] mux_1236_nl;
  wire[0:0] nor_564_nl;
  wire[0:0] nor_565_nl;
  wire[0:0] nor_567_nl;
  wire[0:0] mux_907_nl;
  wire[0:0] or_1393_nl;
  wire[0:0] nor_215_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_194_nl;
  wire[0:0] MultLoop_and_215_nl;
  wire[0:0] MultLoop_and_216_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_136_nl;
  wire[0:0] mux_908_nl;
  wire[0:0] or_1392_nl;
  wire[0:0] nor_214_nl;
  wire[0:0] and_555_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_195_nl;
  wire[0:0] MultLoop_and_212_nl;
  wire[0:0] nor_554_nl;
  wire[0:0] mux_1242_nl;
  wire[0:0] nor_555_nl;
  wire[0:0] nor_556_nl;
  wire[0:0] mux_1244_nl;
  wire[0:0] and_2623_nl;
  wire[0:0] nor_557_nl;
  wire[0:0] and_557_nl;
  wire[0:0] and_560_nl;
  wire[0:0] and_562_nl;
  wire[0:0] mux_919_nl;
  wire[0:0] mux_917_nl;
  wire[0:0] mux_916_nl;
  wire[0:0] or_1358_nl;
  wire[0:0] and_564_nl;
  wire[0:0] mux_923_nl;
  wire[0:0] mux_922_nl;
  wire[0:0] mux_921_nl;
  wire[0:0] mux_920_nl;
  wire[0:0] mux_927_nl;
  wire[0:0] and_571_nl;
  wire[0:0] and_574_nl;
  wire[0:0] mux_929_nl;
  wire[0:0] and_577_nl;
  wire[0:0] and_580_nl;
  wire[0:0] mux_931_nl;
  wire[0:0] and_583_nl;
  wire[0:0] and_585_nl;
  wire[0:0] mux_932_nl;
  wire[0:0] and_610_nl;
  wire[0:0] mux_938_nl;
  wire[0:0] and_624_nl;
  wire[0:0] mux_800_nl;
  wire[0:0] and_727_nl;
  wire[0:0] mux_1247_nl;
  wire[0:0] or_1868_nl;
  wire[0:0] or_1867_nl;
  wire[0:0] ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_nor_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_368_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_183_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_1_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_366_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_182_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_2_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_364_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_181_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_3_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_362_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_180_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_4_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_360_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_179_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_5_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_358_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_178_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_6_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_356_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_177_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_7_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_354_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_176_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_8_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_352_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_175_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_9_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_350_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_174_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_10_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_348_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_173_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_11_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_346_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_172_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_12_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_344_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_171_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_13_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_342_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_170_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_14_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_340_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_169_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_15_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_338_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_168_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_16_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_336_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_167_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_17_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_334_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_166_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_18_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_332_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_165_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_19_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_330_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_164_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_20_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_328_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_163_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_21_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_326_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_162_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_22_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_324_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_161_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_23_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_322_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_160_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_24_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_320_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_159_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_25_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_318_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_158_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_26_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_316_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_157_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_27_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_314_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_156_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_28_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_312_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_155_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_29_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_310_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_154_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_30_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_308_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_153_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_31_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_306_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_152_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_32_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_304_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_151_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_33_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_302_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_150_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_34_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_300_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_149_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_35_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_298_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_148_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_36_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_296_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_147_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_37_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_294_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_146_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_38_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_292_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_145_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_39_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_290_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_144_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_40_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_288_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_143_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_41_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_286_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_142_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_42_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_284_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_141_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_43_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_282_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_140_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_44_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_280_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_139_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_45_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_278_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_138_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_46_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_276_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_137_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_47_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_274_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_136_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_48_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_272_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_135_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_49_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_270_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_134_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_50_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_268_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_133_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_51_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_266_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_132_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_52_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_264_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_131_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_53_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_262_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_130_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_54_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_260_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_129_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_55_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_258_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_128_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_56_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_256_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_127_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_57_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_254_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_126_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_58_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_252_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_125_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_59_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_250_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_124_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_60_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_248_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_123_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_61_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_246_nl;
  wire[0:0] nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_122_nl;
  wire[14:0] IndexLoop_ir_mux_nl;
  wire[14:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_2_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl;
  wire[14:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_2_nor_2_nl;
  wire[0:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_2_and_nl;
  wire[0:0] nor_373_nl;
  wire[0:0] mux_884_nl;
  wire[0:0] or_12_nl;
  wire[0:0] or_1283_nl;
  wire[6:0] IndexLoop_acc_nl;
  wire[7:0] nl_IndexLoop_acc_nl;
  wire[6:0] ReuseLoop_acc_nl;
  wire[7:0] nl_ReuseLoop_acc_nl;
  wire[5:0] IndexLoop_if_acc_13_nl;
  wire[6:0] nl_IndexLoop_if_acc_13_nl;
  wire[6:0] IndexLoop_if_acc_10_nl;
  wire[7:0] nl_IndexLoop_if_acc_10_nl;
  wire[1:0] IndexLoop_if_acc_15_nl;
  wire[2:0] nl_IndexLoop_if_acc_15_nl;
  wire[7:0] IndexLoop_if_acc_8_nl;
  wire[10:0] nl_IndexLoop_if_acc_8_nl;
  wire[3:0] IndexLoop_if_acc_12_nl;
  wire[5:0] nl_IndexLoop_if_acc_12_nl;
  wire[14:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_1_nor_2_nl;
  wire[0:0] nnet_softmax_layer6_t_result_t_softmax_config7_for_1_and_nl;
  wire[0:0] or_1409_nl;
  wire[0:0] or_609_nl;
  wire[0:0] mux_479_nl;
  wire[0:0] mux_487_nl;
  wire[0:0] mux_512_nl;
  wire[0:0] mux_540_nl;
  wire[0:0] mux_542_nl;
  wire[0:0] mux_585_nl;
  wire[0:0] mux_609_nl;
  wire[0:0] mux_453_nl;
  wire[0:0] or_1391_nl;
  wire[0:0] mux_924_nl;
  wire[0:0] mux_499_nl;
  wire[0:0] mux_563_nl;
  wire[0:0] mux_568_nl;
  wire[0:0] mux_579_nl;
  wire[0:0] mux_582_nl;
  wire[0:0] mux_761_nl;
  wire[0:0] mux_4_nl;
  wire[0:0] mux_3_nl;
  wire[0:0] mux_1_nl;
  wire[0:0] mux_762_nl;
  wire[0:0] or_867_nl;
  wire[0:0] mux_481_nl;
  wire[0:0] mux_764_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] or_11_nl;
  wire[0:0] mux_988_nl;
  wire[0:0] nor_450_nl;
  wire[0:0] mux_966_nl;
  wire[0:0] mux_967_nl;
  wire[0:0] nor_441_nl;
  wire[0:0] mux_968_nl;
  wire[0:0] nor_439_nl;
  wire[0:0] nor_440_nl;
  wire[0:0] mux_969_nl;
  wire[0:0] nor_437_nl;
  wire[0:0] nor_438_nl;
  wire[0:0] mux_970_nl;
  wire[0:0] nor_435_nl;
  wire[0:0] nor_436_nl;
  wire[0:0] mux_971_nl;
  wire[0:0] nor_434_nl;
  wire[0:0] mux_972_nl;
  wire[0:0] nor_432_nl;
  wire[0:0] nor_433_nl;
  wire[0:0] mux_973_nl;
  wire[0:0] nor_430_nl;
  wire[0:0] nor_431_nl;
  wire[0:0] mux_974_nl;
  wire[0:0] nor_428_nl;
  wire[0:0] nor_429_nl;
  wire[0:0] mux_975_nl;
  wire[0:0] mux_976_nl;
  wire[0:0] nor_425_nl;
  wire[0:0] nor_426_nl;
  wire[0:0] mux_977_nl;
  wire[0:0] nor_423_nl;
  wire[0:0] nor_424_nl;
  wire[0:0] mux_978_nl;
  wire[0:0] nor_421_nl;
  wire[0:0] nor_422_nl;
  wire[0:0] mux_979_nl;
  wire[0:0] nor_419_nl;
  wire[0:0] nor_420_nl;
  wire[0:0] mux_980_nl;
  wire[0:0] mux_981_nl;
  wire[0:0] nand_150_nl;
  wire[0:0] or_1473_nl;
  wire[0:0] nor_415_nl;
  wire[0:0] nor_416_nl;
  wire[0:0] nor_413_nl;
  wire[0:0] nor_414_nl;
  wire[0:0] mux_984_nl;
  wire[0:0] or_nl;
  wire[0:0] or_1472_nl;
  wire[0:0] mux_985_nl;
  wire[0:0] nor_409_nl;
  wire[0:0] nor_410_nl;
  wire[0:0] mux_986_nl;
  wire[0:0] or_1476_nl;
  wire[0:0] nand_151_nl;
  wire[0:0] mux_987_nl;
  wire[0:0] mux_1095_nl;
  wire[0:0] mux_1094_nl;
  wire[0:0] mux_1093_nl;
  wire[0:0] or_1621_nl;
  wire[0:0] or_1620_nl;
  wire[0:0] or_1619_nl;
  wire[0:0] or_1629_nl;
  wire[0:0] mux_1102_nl;
  wire[0:0] mux_1101_nl;
  wire[0:0] or_1628_nl;
  wire[0:0] mux_1136_nl;
  wire[0:0] mux_1135_nl;
  wire[0:0] mux_1134_nl;
  wire[0:0] nor_629_nl;
  wire[0:0] nor_630_nl;
  wire[0:0] nor_631_nl;
  wire[0:0] nor_632_nl;
  wire[0:0] mux_1195_nl;
  wire[0:0] nor_577_nl;
  wire[0:0] mux_1209_nl;
  wire[0:0] nor_574_nl;
  wire[0:0] nor_575_nl;
  wire[0:0] mux_1214_nl;
  wire[0:0] or_1819_nl;
  wire[0:0] or_1818_nl;
  wire[0:0] or_1823_nl;
  wire[0:0] or_1822_nl;
  wire[0:0] ReuseLoop_mux1h_3_nl;
  wire[7:0] acc_nl;
  wire[8:0] nl_acc_nl;
  wire[5:0] ReuseLoop_1_ReuseLoop_1_mux_1_nl;
  wire[0:0] ReuseLoop_1_or_3_nl;
  wire[0:0] ReuseLoop_1_or_4_nl;
  wire[3:0] ReuseLoop_2_acc_nl;
  wire[4:0] nl_ReuseLoop_2_acc_nl;
  wire[2:0] ReuseLoop_2_mux_1_nl;
  wire[0:0] and_2668_nl;
  wire[0:0] ac_math_ac_reciprocal_pwl_AC_TRN_71_51_false_AC_TRN_AC_WRAP_91_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_71_51_false_AC_TRN_AC_WRAP_91_21_false_AC_TRN_AC_WRAP_output_pwl_or_1_nl;
  wire[9:0] ac_math_ac_reciprocal_pwl_AC_TRN_71_51_false_AC_TRN_AC_WRAP_91_21_false_AC_TRN_AC_WRAP_output_pwl_mux1h_2_nl;
  wire[8:0] ac_math_ac_reciprocal_pwl_AC_TRN_71_51_false_AC_TRN_AC_WRAP_91_21_false_AC_TRN_AC_WRAP_output_pwl_mux1h_3_nl;
  wire[5:0] ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_qif_mux_2_nl;
  wire[0:0] ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_qif_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_qif_and_1_nl;
  wire[0:0] ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_qif_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_qif_or_1_nl;
  wire[0:0] SUM_EXP_LOOP_SUM_EXP_LOOP_and_5_nl;
  wire[0:0] SUM_EXP_LOOP_SUM_EXP_LOOP_and_6_nl;
  wire[0:0] SUM_EXP_LOOP_mux_3_nl;
  wire[67:0] SUM_EXP_LOOP_SUM_EXP_LOOP_mux_2_nl;
  wire[0:0] SUM_EXP_LOOP_or_1_nl;
  wire[0:0] SUM_EXP_LOOP_SUM_EXP_LOOP_and_7_nl;
  wire[67:0] SUM_EXP_LOOP_mux1h_5_nl;
  wire[8:0] ReuseLoop_if_mux_2_nl;
  wire[0:0] ReuseLoop_and_4_nl;
  wire[0:0] ReuseLoop_mux1h_5_nl;
  wire[14:0] ReuseLoop_and_5_nl;
  wire[14:0] ReuseLoop_mux1h_6_nl;
  wire[7:0] ReuseLoop_ReuseLoop_and_2_nl;
  wire[7:0] ReuseLoop_mux_1_nl;
  wire[0:0] not_3912_nl;
  wire[10:0] ReuseLoop_ReuseLoop_mux_1_nl;
  wire[0:0] IndexLoop_if_mux1h_5_nl;
  wire[14:0] IndexLoop_if_mux1h_6_nl;
  wire[0:0] IndexLoop_if_mux1h_7_nl;
  wire[0:0] IndexLoop_if_mux1h_8_nl;
  wire[0:0] IndexLoop_if_IndexLoop_if_and_2_nl;
  wire[0:0] IndexLoop_if_IndexLoop_if_and_3_nl;
  wire[0:0] IndexLoop_if_IndexLoop_if_or_1_nl;
  wire[17:0] IndexLoop_if_IndexLoop_if_mux_1_nl;
  wire[17:0] ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_80_nl;
  wire[18:0] nl_ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_80_nl;
  wire[0:0] ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_17_nl;
  wire[14:0] ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_18_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_mux_2_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_mux_3_nl;
  wire[157:0] mul_1_nl;
  wire signed [159:0] nl_mul_1_nl;
  wire[66:0] nnet_product_input_t_config2_weight_t_config2_accum_t_1_mux1h_3_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_1_or_2_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_1_nnet_product_input_t_config2_weight_t_config2_accum_t_1_and_1_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_1_mux_3_nl;
  wire[73:0] nnet_product_input_t_config2_weight_t_config2_accum_t_1_mux1h_4_nl;
  wire[16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_1_mux1h_5_nl;
  wire[27:0] mul_2_nl;
  wire signed [35:0] nl_mul_2_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_1_mux_4_nl;
  wire[17:0] MultLoop_mux_325_nl;
  wire[17:0] MultLoop_mux_326_nl;
  wire[17:0] MultLoop_mux_327_nl;
  wire[17:0] MultLoop_mux_328_nl;
  wire[17:0] MultLoop_mux_329_nl;
  wire[17:0] MultLoop_mux_330_nl;
  wire[17:0] MultLoop_mux_331_nl;
  wire[17:0] MultLoop_mux_332_nl;
  wire[17:0] MultLoop_mux_333_nl;
  wire[17:0] MultLoop_mux_334_nl;
  wire[17:0] MultLoop_mux_335_nl;
  wire[17:0] MultLoop_mux_336_nl;
  wire[17:0] MultLoop_mux_337_nl;
  wire[17:0] MultLoop_mux_338_nl;
  wire[17:0] MultLoop_mux_339_nl;
  wire[17:0] MultLoop_mux_340_nl;
  wire[17:0] MultLoop_mux_341_nl;
  wire[17:0] MultLoop_mux_342_nl;
  wire[17:0] MultLoop_mux_343_nl;
  wire[17:0] MultLoop_mux_344_nl;
  wire[17:0] MultLoop_mux_345_nl;
  wire[17:0] MultLoop_mux_346_nl;
  wire[17:0] MultLoop_mux_347_nl;
  wire[17:0] MultLoop_mux_348_nl;
  wire[17:0] MultLoop_mux_349_nl;
  wire[17:0] MultLoop_mux_350_nl;
  wire[17:0] MultLoop_mux_351_nl;
  wire[17:0] MultLoop_mux_352_nl;
  wire[17:0] MultLoop_mux_353_nl;
  wire[17:0] MultLoop_mux_354_nl;
  wire[17:0] MultLoop_mux_355_nl;
  wire[17:0] MultLoop_mux_356_nl;
  wire[17:0] MultLoop_mux_357_nl;
  wire[17:0] MultLoop_mux_358_nl;
  wire[17:0] MultLoop_mux_359_nl;
  wire[17:0] MultLoop_mux_360_nl;
  wire[17:0] MultLoop_mux_361_nl;
  wire[17:0] MultLoop_mux_362_nl;
  wire[17:0] MultLoop_mux_363_nl;
  wire[17:0] MultLoop_mux_364_nl;
  wire[17:0] MultLoop_mux_365_nl;
  wire[17:0] MultLoop_mux_366_nl;
  wire[17:0] MultLoop_mux_367_nl;
  wire[17:0] MultLoop_mux_368_nl;
  wire[17:0] MultLoop_mux_369_nl;
  wire[17:0] MultLoop_mux_370_nl;
  wire[17:0] MultLoop_mux_371_nl;
  wire[17:0] MultLoop_mux_372_nl;
  wire[17:0] MultLoop_mux_373_nl;
  wire[17:0] MultLoop_mux_374_nl;
  wire[17:0] MultLoop_mux_375_nl;
  wire[17:0] MultLoop_mux_376_nl;
  wire[17:0] MultLoop_mux_377_nl;
  wire[17:0] MultLoop_mux_378_nl;
  wire[17:0] MultLoop_mux_379_nl;
  wire[17:0] MultLoop_mux_380_nl;
  wire[17:0] MultLoop_mux_381_nl;
  wire[17:0] MultLoop_mux_382_nl;
  wire[17:0] MultLoop_mux_383_nl;
  wire[17:0] MultLoop_mux_384_nl;
  wire[17:0] MultLoop_mux_385_nl;
  wire[17:0] MultLoop_mux_386_nl;
  wire[17:0] MultLoop_mux_387_nl;
  wire[17:0] MultLoop_mux_388_nl;
  wire[17:0] MultLoop_mux_389_nl;
  wire[17:0] MultLoop_mux_390_nl;
  wire[0:0] MultLoop_or_9_nl;
  wire[17:0] MultLoop_mux1h_66_nl;
  wire[27:0] MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_1_nl;
  wire signed [35:0] nl_MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_1_nl;
  wire[17:0] MultLoop_mux1h_67_nl;
  wire[22:0] operator_18_8_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_operator_18_8_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[0:0] operator_18_8_true_AC_TRN_AC_WRAP_1_mux1h_5_nl;
  wire[3:0] operator_18_8_true_AC_TRN_AC_WRAP_1_mux1h_6_nl;
  wire[12:0] operator_18_8_true_AC_TRN_AC_WRAP_1_mux1h_7_nl;
  wire[3:0] operator_18_8_true_AC_TRN_AC_WRAP_1_nor_1_nl;
  wire[3:0] operator_18_8_true_AC_TRN_AC_WRAP_1_mux1h_8_nl;
  wire[18:0] operator_18_8_true_AC_TRN_AC_WRAP_1_operator_18_8_true_AC_TRN_AC_WRAP_1_operator_18_8_true_AC_TRN_AC_WRAP_1_and_nl;
  wire[18:0] ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_79_nl;
  wire[19:0] nl_ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_79_nl;
  wire[1:0] operator_18_8_true_AC_TRN_AC_WRAP_1_operator_18_8_true_AC_TRN_AC_WRAP_1_mux_1_nl;
  wire[0:0] SUM_EXP_LOOP_SUM_EXP_LOOP_and_8_nl;
  wire[66:0] SUM_EXP_LOOP_mux1h_6_nl;
  wire[0:0] SUM_EXP_LOOP_SUM_EXP_LOOP_and_9_nl;
  wire[66:0] SUM_EXP_LOOP_mux1h_7_nl;
  wire[4:0] mux_1250_nl;
  wire[2:0] mux_1249_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [2:0] nl_U_ROM_1i3_1o10_bb905e8578f158e8f5b59add1dc96bdb2f_rg_I_1;
  assign nl_U_ROM_1i3_1o10_bb905e8578f158e8f5b59add1dc96bdb2f_rg_I_1 = operator_71_0_false_AC_TRN_AC_WRAP_lshift_itm[69:67];
  wire [70:0] nl_operator_91_21_false_AC_TRN_AC_WRAP_rshift_rg_a;
  assign nl_operator_91_21_false_AC_TRN_AC_WRAP_rshift_rg_a = {z_out_2 , (z_out_17[9:0])
      , 50'b00000000000000000000000000000000000000000000000000};
  wire [7:0] nl_operator_91_21_false_AC_TRN_AC_WRAP_rshift_rg_s;
  assign nl_operator_91_21_false_AC_TRN_AC_WRAP_rshift_rg_s = {z_out_3 , (~ (libraries_leading_sign_71_0_e5d4bd9dc928fda5adf5bf26ec9a2550b9a2_1[1:0]))};
  wire [8:0] nl_U_ROM_1i9_1o3_2fa806bf16b3e0d54016201674d036b62f_rg_I_1;
  assign nl_U_ROM_1i9_1o3_2fa806bf16b3e0d54016201674d036b62f_rg_I_1 = reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2[8:0];
  wire [2:0] nl_U_ROM_1i3_1o8_bdb5a3eca137308489a677a1241b230a2e_rg_I_1;
  assign nl_U_ROM_1i3_1o8_bdb5a3eca137308489a677a1241b230a2e_rg_I_1 = operator_71_0_false_AC_TRN_AC_WRAP_lshift_itm[69:67];
  wire [69:0] nl_operator_71_0_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_operator_71_0_false_AC_TRN_AC_WRAP_lshift_rg_a = z_out_10[69:0];
  wire [70:0] nl_leading_sign_71_0_rg_mantissa;
  assign nl_leading_sign_71_0_rg_mantissa = z_out_10;
  wire[10:0] ac_math_ac_pow2_pwl_AC_TRN_19_7_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_ac_math_ac_pow2_pwl_AC_TRN_19_7_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[2:0] mux_1248_nl;
  wire[6:0] mux_1251_nl;
  wire [20:0] nl_CALC_EXP_LOOP_10_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign mux_1248_nl = MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, z_out_12[12:11]);
  assign mux_1251_nl = MUX_v_7_4_2(7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111,
      z_out_12[12:11]);
  assign nl_ac_math_ac_pow2_pwl_AC_TRN_19_7_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = ({(mux_1248_nl) , 1'b1 , (mux_1251_nl)}) + conv_u2u_9_11(z_out_25[18:10]);
  assign ac_math_ac_pow2_pwl_AC_TRN_19_7_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_ac_math_ac_pow2_pwl_AC_TRN_19_7_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_CALC_EXP_LOOP_10_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_a = {(ac_math_ac_pow2_pwl_AC_TRN_19_7_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl)
      , (z_out_25[9:0])};
  wire [6:0] nl_CALC_EXP_LOOP_10_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_CALC_EXP_LOOP_10_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_s = z_out_12[19:13];
  wire [179:0] nl_mnist_mlp_core_layer7_out_rsci_inst_layer7_out_rsci_idat;
  assign nl_mnist_mlp_core_layer7_out_rsci_inst_layer7_out_rsci_idat = {6'b000000
      , layer7_out_rsci_idat_173_162 , 6'b000000 , layer7_out_rsci_idat_155_144 ,
      6'b000000 , layer7_out_rsci_idat_137_126 , 6'b000000 , layer7_out_rsci_idat_119_108
      , 6'b000000 , layer7_out_rsci_idat_101_90 , 6'b000000 , layer7_out_rsci_idat_83_72
      , 6'b000000 , layer7_out_rsci_idat_65_54 , 6'b000000 , layer7_out_rsci_idat_47_36
      , 6'b000000 , layer7_out_rsci_idat_29_18 , 6'b000000 , layer7_out_rsci_idat_11_0};
  wire [1:0] nl_mnist_mlp_core_w2_rsci_1_inst_w2_rsci_adra_d_core_psct;
  assign nl_mnist_mlp_core_w2_rsci_1_inst_w2_rsci_adra_d_core_psct = {and_dcpl_82
      , and_dcpl_82};
  wire [1:0] nl_mnist_mlp_core_w2_rsci_1_inst_w2_rsci_ena_d_core_psct;
  assign nl_mnist_mlp_core_w2_rsci_1_inst_w2_rsci_ena_d_core_psct = {and_dcpl_82
      , and_dcpl_82};
  wire [1:0] nl_mnist_mlp_core_w2_rsci_1_inst_w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_mnist_mlp_core_w2_rsci_1_inst_w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = {and_dcpl_82 , and_dcpl_82};
  wire[6:0] MultLoop_1_acc_1_nl;
  wire[7:0] nl_MultLoop_1_acc_1_nl;
  wire [31:0] nl_mnist_mlp_core_w2_rsci_1_inst_w2_rsci_adra_d_core_pff;
  assign nl_MultLoop_1_acc_1_nl = conv_u2u_6_7({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_2_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_4_reg
      , (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2[10:9])})
      + 7'b0110001;
  assign MultLoop_1_acc_1_nl = nl_MultLoop_1_acc_1_nl[6:0];
  assign nl_mnist_mlp_core_w2_rsci_1_inst_w2_rsci_adra_d_core_pff = {(MultLoop_1_acc_1_nl)
      , (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2[8:0])
      , 1'b0 , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_2_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_4_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2};
  wire [1:0] nl_mnist_mlp_core_w4_rsci_1_inst_w4_rsci_ena_d_core_psct;
  assign nl_mnist_mlp_core_w4_rsci_1_inst_w4_rsci_ena_d_core_psct = {and_dcpl_77
      , and_dcpl_77};
  wire [1:0] nl_mnist_mlp_core_w4_rsci_1_inst_w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_mnist_mlp_core_w4_rsci_1_inst_w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = {and_dcpl_77 , and_dcpl_77};
  wire [1:0] nl_mnist_mlp_core_w4_rsci_1_inst_w4_rsci_adra_d_core_psct_pff;
  assign nl_mnist_mlp_core_w4_rsci_1_inst_w4_rsci_adra_d_core_psct_pff = {and_dcpl_77
      , and_dcpl_77};
  wire [23:0] nl_mnist_mlp_core_w4_rsci_1_inst_w4_rsci_adra_d_core_pff;
  assign nl_mnist_mlp_core_w4_rsci_1_inst_w4_rsci_adra_d_core_pff = {1'b1 , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2
      , 1'b0 , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2};
  wire [1:0] nl_mnist_mlp_core_w6_rsci_1_inst_w6_rsci_adra_d_core_psct;
  assign nl_mnist_mlp_core_w6_rsci_1_inst_w6_rsci_adra_d_core_psct = {and_73_rmff
      , and_73_rmff};
  wire [1:0] nl_mnist_mlp_core_w6_rsci_1_inst_w6_rsci_ena_d_core_psct;
  assign nl_mnist_mlp_core_w6_rsci_1_inst_w6_rsci_ena_d_core_psct = {and_73_rmff
      , and_73_rmff};
  wire [1:0] nl_mnist_mlp_core_w6_rsci_1_inst_w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_mnist_mlp_core_w6_rsci_1_inst_w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = {and_73_rmff , and_73_rmff};
  wire [19:0] nl_mnist_mlp_core_w6_rsci_1_inst_w6_rsci_adra_d_core_pff;
  assign nl_mnist_mlp_core_w6_rsci_1_inst_w6_rsci_adra_d_core_pff = {(z_out_2[3:0])
      , (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2[5:0])
      , 1'b0 , (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2[8:0])};
  wire [0:0] nl_mnist_mlp_core_core_fsm_inst_InitAccumLoop_C_0_tr0;
  assign nl_mnist_mlp_core_core_fsm_inst_InitAccumLoop_C_0_tr0 = z_out[6];
  wire [0:0] nl_mnist_mlp_core_core_fsm_inst_IndexLoop_C_0_tr0;
  assign nl_mnist_mlp_core_core_fsm_inst_IndexLoop_C_0_tr0 = ~ IndexLoop_stage_0;
  wire [0:0] nl_mnist_mlp_core_core_fsm_inst_InitAccumLoop_1_C_0_tr0;
  assign nl_mnist_mlp_core_core_fsm_inst_InitAccumLoop_1_C_0_tr0 = z_out[6];
  wire [0:0] nl_mnist_mlp_core_core_fsm_inst_ReuseLoop_1_C_0_tr0;
  assign nl_mnist_mlp_core_core_fsm_inst_ReuseLoop_1_C_0_tr0 = ~ IndexLoop_stage_0;
  wire [0:0] nl_mnist_mlp_core_core_fsm_inst_InitAccumLoop_2_C_0_tr0;
  assign nl_mnist_mlp_core_core_fsm_inst_InitAccumLoop_2_C_0_tr0 = ~ z_out_1_3;
  wire [0:0] nl_mnist_mlp_core_core_fsm_inst_ReuseLoop_2_C_0_tr0;
  assign nl_mnist_mlp_core_core_fsm_inst_ReuseLoop_2_C_0_tr0 = ~ IndexLoop_stage_0;
  wire [0:0] nl_mnist_mlp_core_core_fsm_inst_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_C_0_tr0;
  assign nl_mnist_mlp_core_core_fsm_inst_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_C_0_tr0
      = ~ IndexLoop_stage_0;
  ccs_in_v1 #(.rscid(32'sd6),
  .width(32'sd1152)) b2_rsci (
      .dat(b2_rsc_dat),
      .idat(b2_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd8),
  .width(32'sd1152)) b4_rsci (
      .dat(b4_rsc_dat),
      .idat(b4_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd10),
  .width(32'sd180)) b6_rsci (
      .dat(b6_rsc_dat),
      .idat(b6_rsci_idat)
    );
  ROM_1i3_1o10_2c1f806487d17904bea969f4e53173bcb1  U_ROM_1i3_1o10_bb905e8578f158e8f5b59add1dc96bdb2f_rg
      (
      .I_1(nl_U_ROM_1i3_1o10_bb905e8578f158e8f5b59add1dc96bdb2f_rg_I_1[2:0]),
      .O_1(ROM_1i3_1o10_bb905e8578f158e8f5b59add1dc96bdb2f_1)
    );
  mgc_shift_br_v5 #(.width_a(32'sd71),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd91)) operator_91_21_false_AC_TRN_AC_WRAP_rshift_rg (
      .a(nl_operator_91_21_false_AC_TRN_AC_WRAP_rshift_rg_a[70:0]),
      .s(nl_operator_91_21_false_AC_TRN_AC_WRAP_rshift_rg_s[7:0]),
      .z(operator_91_21_false_AC_TRN_AC_WRAP_rshift_itm)
    );
  ROM_1i11_1o5_35e12f400da6925eda56234f89e8055db3  U_ROM_1i11_1o5_b94ddd86102738ded3ce1c444a799cda31_rg
      (
      .I_1(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2),
      .O_1(ROM_1i11_1o5_b94ddd86102738ded3ce1c444a799cda31_1)
    );
  ROM_1i9_1o3_0cffcd7ae8128c5cac71e8022405e1ebb1  U_ROM_1i9_1o3_2fa806bf16b3e0d54016201674d036b62f_rg
      (
      .I_1(nl_U_ROM_1i9_1o3_2fa806bf16b3e0d54016201674d036b62f_rg_I_1[8:0]),
      .O_1(ROM_1i9_1o3_2fa806bf16b3e0d54016201674d036b62f_1)
    );
  ROM_1i3_1o8_b7f1baaf117249900fa3606aa9bde444b0  U_ROM_1i3_1o8_bdb5a3eca137308489a677a1241b230a2e_rg
      (
      .I_1(nl_U_ROM_1i3_1o8_bdb5a3eca137308489a677a1241b230a2e_rg_I_1[2:0]),
      .O_1(ROM_1i3_1o8_bdb5a3eca137308489a677a1241b230a2e_1)
    );
  mgc_shift_l_v5 #(.width_a(32'sd70),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd70)) operator_71_0_false_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_operator_71_0_false_AC_TRN_AC_WRAP_lshift_rg_a[69:0]),
      .s(libraries_leading_sign_71_0_e5d4bd9dc928fda5adf5bf26ec9a2550b9a2_1),
      .z(operator_71_0_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  leading_sign_71_0  leading_sign_71_0_rg (
      .mantissa(nl_leading_sign_71_0_rg_mantissa[70:0]),
      .rtn(libraries_leading_sign_71_0_e5d4bd9dc928fda5adf5bf26ec9a2550b9a2_1)
    );
  mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd67)) CALC_EXP_LOOP_10_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(nl_CALC_EXP_LOOP_10_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(nl_CALC_EXP_LOOP_10_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_s[6:0]),
      .z(z_out_9)
    );
  mnist_mlp_core_input1_rsci mnist_mlp_core_input1_rsci_inst (
      .clk(clk),
      .rst(rst),
      .input1_rsc_dat(input1_rsc_dat),
      .input1_rsc_vld(input1_rsc_vld),
      .input1_rsc_rdy(input1_rsc_rdy),
      .core_wen(core_wen),
      .input1_rsci_oswt(reg_w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_0_cse),
      .input1_rsci_wen_comp(input1_rsci_wen_comp),
      .input1_rsci_idat_mxwt(input1_rsci_idat_mxwt)
    );
  mnist_mlp_core_layer7_out_rsci mnist_mlp_core_layer7_out_rsci_inst (
      .clk(clk),
      .rst(rst),
      .layer7_out_rsc_dat(layer7_out_rsc_dat),
      .layer7_out_rsc_vld(layer7_out_rsc_vld),
      .layer7_out_rsc_rdy(layer7_out_rsc_rdy),
      .core_wen(core_wen),
      .layer7_out_rsci_oswt(reg_layer7_out_rsci_ivld_core_psct_cse),
      .layer7_out_rsci_wen_comp(layer7_out_rsci_wen_comp),
      .layer7_out_rsci_idat(nl_mnist_mlp_core_layer7_out_rsci_inst_layer7_out_rsci_idat[179:0])
    );
  mnist_mlp_core_const_size_in_1_rsci mnist_mlp_core_const_size_in_1_rsci_inst (
      .clk(clk),
      .rst(rst),
      .const_size_in_1_rsc_dat(const_size_in_1_rsc_dat),
      .const_size_in_1_rsc_vld(const_size_in_1_rsc_vld),
      .const_size_in_1_rsc_rdy(const_size_in_1_rsc_rdy),
      .core_wen(core_wen),
      .const_size_in_1_rsci_oswt(reg_const_size_out_1_rsci_ivld_core_psct_cse),
      .const_size_in_1_rsci_wen_comp(const_size_in_1_rsci_wen_comp)
    );
  mnist_mlp_core_const_size_out_1_rsci mnist_mlp_core_const_size_out_1_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .const_size_out_1_rsc_dat(const_size_out_1_rsc_dat),
      .const_size_out_1_rsc_vld(const_size_out_1_rsc_vld),
      .const_size_out_1_rsc_rdy(const_size_out_1_rsc_rdy),
      .core_wen(core_wen),
      .const_size_out_1_rsci_oswt(reg_const_size_out_1_rsci_ivld_core_psct_cse),
      .const_size_out_1_rsci_wen_comp(const_size_out_1_rsci_wen_comp)
    );
  mnist_mlp_core_w2_rsci_1 mnist_mlp_core_w2_rsci_1_inst (
      .clk(clk),
      .rst(rst),
      .w2_rsci_adra_d(w2_rsci_adra_d_reg),
      .w2_rsci_ena_d(w2_rsci_ena_d_reg),
      .w2_rsci_qa_d(w2_rsci_qa_d),
      .w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .w2_rsci_oswt(reg_w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_0_cse),
      .w2_rsci_adra_d_core_psct(nl_mnist_mlp_core_w2_rsci_1_inst_w2_rsci_adra_d_core_psct[1:0]),
      .w2_rsci_ena_d_core_psct(nl_mnist_mlp_core_w2_rsci_1_inst_w2_rsci_ena_d_core_psct[1:0]),
      .w2_rsci_qa_d_mxwt(w2_rsci_qa_d_mxwt),
      .w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_mnist_mlp_core_w2_rsci_1_inst_w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[1:0]),
      .w2_rsci_adra_d_core_pff(nl_mnist_mlp_core_w2_rsci_1_inst_w2_rsci_adra_d_core_pff[31:0]),
      .w2_rsci_oswt_pff(and_dcpl_82)
    );
  mnist_mlp_core_w4_rsci_1 mnist_mlp_core_w4_rsci_1_inst (
      .clk(clk),
      .rst(rst),
      .w4_rsci_adra_d(w4_rsci_adra_d_reg),
      .w4_rsci_ena_d(w4_rsci_ena_d_reg),
      .w4_rsci_qa_d(w4_rsci_qa_d),
      .w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .w4_rsci_oswt(reg_w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_0_cse),
      .w4_rsci_ena_d_core_psct(nl_mnist_mlp_core_w4_rsci_1_inst_w4_rsci_ena_d_core_psct[1:0]),
      .w4_rsci_qa_d_mxwt(w4_rsci_qa_d_mxwt),
      .w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_mnist_mlp_core_w4_rsci_1_inst_w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[1:0]),
      .w4_rsci_adra_d_core_psct_pff(nl_mnist_mlp_core_w4_rsci_1_inst_w4_rsci_adra_d_core_psct_pff[1:0]),
      .w4_rsci_oswt_pff(and_dcpl_77),
      .w4_rsci_adra_d_core_pff(nl_mnist_mlp_core_w4_rsci_1_inst_w4_rsci_adra_d_core_pff[23:0])
    );
  mnist_mlp_core_w6_rsci_1 mnist_mlp_core_w6_rsci_1_inst (
      .clk(clk),
      .rst(rst),
      .w6_rsci_adra_d(w6_rsci_adra_d_reg),
      .w6_rsci_ena_d(w6_rsci_ena_d_reg),
      .w6_rsci_qa_d(w6_rsci_qa_d),
      .w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .w6_rsci_oswt(reg_w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_0_cse),
      .w6_rsci_adra_d_core_psct(nl_mnist_mlp_core_w6_rsci_1_inst_w6_rsci_adra_d_core_psct[1:0]),
      .w6_rsci_ena_d_core_psct(nl_mnist_mlp_core_w6_rsci_1_inst_w6_rsci_ena_d_core_psct[1:0]),
      .w6_rsci_qa_d_mxwt(w6_rsci_qa_d_mxwt),
      .w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_mnist_mlp_core_w6_rsci_1_inst_w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[1:0]),
      .w6_rsci_adra_d_core_pff(nl_mnist_mlp_core_w6_rsci_1_inst_w6_rsci_adra_d_core_pff[19:0]),
      .w6_rsci_oswt_pff(and_73_rmff)
    );
  mnist_mlp_core_staller mnist_mlp_core_staller_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .input1_rsci_wen_comp(input1_rsci_wen_comp),
      .layer7_out_rsci_wen_comp(layer7_out_rsci_wen_comp),
      .const_size_in_1_rsci_wen_comp(const_size_in_1_rsci_wen_comp),
      .const_size_out_1_rsci_wen_comp(const_size_out_1_rsci_wen_comp)
    );
  mnist_mlp_core_core_fsm mnist_mlp_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output),
      .InitAccumLoop_C_0_tr0(nl_mnist_mlp_core_core_fsm_inst_InitAccumLoop_C_0_tr0[0:0]),
      .IndexLoop_C_0_tr0(nl_mnist_mlp_core_core_fsm_inst_IndexLoop_C_0_tr0[0:0]),
      .InitAccumLoop_1_C_0_tr0(nl_mnist_mlp_core_core_fsm_inst_InitAccumLoop_1_C_0_tr0[0:0]),
      .ReuseLoop_1_C_0_tr0(nl_mnist_mlp_core_core_fsm_inst_ReuseLoop_1_C_0_tr0[0:0]),
      .InitAccumLoop_2_C_0_tr0(nl_mnist_mlp_core_core_fsm_inst_InitAccumLoop_2_C_0_tr0[0:0]),
      .ReuseLoop_2_C_0_tr0(nl_mnist_mlp_core_core_fsm_inst_ReuseLoop_2_C_0_tr0[0:0]),
      .nnet_softmax_layer6_t_result_t_softmax_config7_for_1_C_0_tr0(nl_mnist_mlp_core_core_fsm_inst_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_C_0_tr0[0:0])
    );
  assign and_73_rmff = and_dcpl_70 & nor_298_cse & and_817_cse & and_dcpl_66;
  assign nor_942_cse = ~((fsm_output[3:2]!=2'b00));
  assign nor_943_cse = ~((fsm_output[5:4]!=2'b00));
  assign nor_944_cse = ~((fsm_output[7:6]!=2'b00));
  assign nor_941_nl = ~(IndexLoop_asn_3_itm_1 | (~ IndexLoop_stage_0_2));
  assign mux_989_cse = MUX_s_1_2_2((InitAccumLoop_1_iacc_6_0_sva_5_0[5]), (nor_941_nl),
      fsm_output[0]);
  assign or_1479_cse = IndexLoop_asn_3_itm_1 | (~ IndexLoop_stage_0_2);
  assign mux_990_cse = MUX_s_1_2_2((InitAccumLoop_1_iacc_6_0_sva_5_0[5]), or_1479_cse,
      fsm_output[0]);
  assign nor_936_cse = ~(mux_990_cse | (InitAccumLoop_1_iacc_6_0_sva_5_0[2]));
  assign nor_937_cse = ~((InitAccumLoop_1_iacc_6_0_sva_5_0[4:3]!=2'b00));
  assign nor_923_cse = ~((InitAccumLoop_1_iacc_6_0_sva_5_0[1:0]!=2'b00));
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse =
      core_wen & (and_dcpl_158 | and_dcpl_60);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_385_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_125_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_383_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_124_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_381_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_123_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_379_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_122_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_377_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_121_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_375_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_120_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_373_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_119_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_371_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_118_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_369_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_117_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_367_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_116_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_365_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_115_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_363_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_114_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_361_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_113_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_359_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_112_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_357_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_111_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_355_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_110_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_353_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_109_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_351_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_108_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_349_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_107_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_347_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_106_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_345_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_105_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_343_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_104_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_341_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_103_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_339_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_102_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_337_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_101_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_335_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_100_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_333_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_99_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_331_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_98_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_329_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_97_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_327_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_96_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_325_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_128_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_263_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_129_cse)
      & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_cse =
      core_wen & (and_dcpl_160 | and_dcpl_55);
  assign nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_15_cse
      = MultLoop_2_MultLoop_2_nor_2_itm_1 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_57_rgt
      = nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_15_cse
      & and_dcpl_55;
  assign nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_14_cse
      = MultLoop_2_and_15_itm_1 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_53_rgt
      = nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_14_cse
      & and_dcpl_55;
  assign nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_13_cse
      = MultLoop_2_and_14_itm_1 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_49_rgt
      = nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_13_cse
      & and_dcpl_55;
  assign nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_or_9_cse =
      or_dcpl_544 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_45_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_or_9_cse)
      & and_dcpl_55;
  assign nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_11_cse
      = MultLoop_2_and_7_itm_1 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_41_rgt
      = nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_11_cse
      & and_dcpl_55;
  assign nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_10_cse
      = MultLoop_2_and_6_itm_1 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_37_rgt
      = nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_10_cse
      & and_dcpl_55;
  assign nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_9_cse
      = MultLoop_2_and_5_itm_1 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_33_rgt
      = nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_9_cse &
      and_dcpl_55;
  assign nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_or_8_cse =
      or_dcpl_540 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_29_rgt
      = (~ nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_or_8_cse)
      & and_dcpl_55;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_and_cse
      = core_wen & (~(or_tmp_91 | (fsm_output[5]) | or_941_cse | (fsm_output[2:0]!=3'b011)
      | (~ IndexLoop_stage_0) | IndexLoop_IndexLoop_nor_tmp));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_1_and_cse = core_wen
      & (~(or_dcpl_469 | or_dcpl_467));
  assign or_381_cse = (~ (fsm_output[2])) | (~ (fsm_output[6])) | (fsm_output[7]);
  assign or_1420_tmp = or_dcpl_539 | (ReuseLoop_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_outidx_const_assign_1_ReuseLoop_2_asn_tmp_3_2_0_psp_sva_1[2]);
  assign and_817_cse = (fsm_output[2:1]==2'b11);
  assign and_810_cse_1 = (fsm_output[1:0]==2'b11);
  assign nor_306_cse = ~((fsm_output[1:0]!=2'b00));
  assign or_864_cse = (fsm_output[7:6]!=2'b10);
  assign or_865_cse_1 = (fsm_output[7:6]!=2'b01);
  assign CALC_SOFTMAX_LOOP_6_or_1_nl = (z_out_18_157_10[147:82]!=66'b000000000000000000000000000000000000000000000000000000000000000000);
  assign CALC_SOFTMAX_LOOP_6_or_cse = MUX_v_12_2_2((z_out_18_157_10[81:70]), 12'b111111111111,
      (CALC_SOFTMAX_LOOP_6_or_1_nl));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_3_and_seb = (reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_reg[5])
      & (~((reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_reg[4:3]==2'b11)));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_3_nor_2_nl = ~(MUX_v_3_2_2((reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_reg[2:0]),
      3'b111, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_3_sva_mx0w1));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_3_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl
      = ~(MUX_v_3_2_2((nnet_softmax_layer6_t_result_t_softmax_config7_for_3_nor_2_nl),
      3'b111, nnet_softmax_layer6_t_result_t_softmax_config7_for_3_and_seb));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_3_nor_3_nl = ~(MUX_v_12_2_2(reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_1_reg,
      12'b111111111111, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_3_sva_mx0w1));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_3_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_1_nl
      = ~(MUX_v_12_2_2((nnet_softmax_layer6_t_result_t_softmax_config7_for_3_nor_3_nl),
      12'b111111111111, nnet_softmax_layer6_t_result_t_softmax_config7_for_3_and_seb));
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_644_nl
      = (~ or_dcpl_490) & and_dcpl_155;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_273_nl =
      (((and_dcpl_181 & and_dcpl_178) | ((~ or_dcpl_447) & and_dcpl_185)) & and_dcpl_65)
      | (and_dcpl_189 & (~ (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[4]))
      & and_dcpl_188 & and_dcpl_60);
  assign or_880_nl = (ReuseLoop_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_outidx_const_assign_1_ReuseLoop_2_asn_tmp_3_2_0_psp_sva_1!=3'b000);
  assign mux_486_nl = MUX_s_1_2_2(and_2658_cse, or_tmp_384, or_880_nl);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_305_nl =
      ((((~ or_dcpl_572) & or_dcpl_447 & and_dcpl_176) | ((~ or_dcpl_572) & or_dcpl_447
      & and_dcpl_185)) & and_dcpl_65) | ((~((or_1420_tmp & and_dcpl_185) | (mux_486_nl)
      | (~ IndexLoop_stage_0_2))) & and_dcpl_55);
  assign and_193_nl = or_dcpl_495 & IndexLoop_stage_0_2 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_652_nl
      = (~(or_dcpl_338 | or_dcpl_344)) & and_dcpl_160;
  assign and_174_nl = and_dcpl_54 & and_dcpl_171 & (~ (fsm_output[1]));
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_192_rgt
      = MUX1HOT_v_18_7_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
      z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_1_sva_1,
      InitAccumLoop_2_slc_InitAccumLoop_2_asn_18_17_0_ctmp_sva_1, ({3'b000 , (nnet_softmax_layer6_t_result_t_softmax_config7_for_3_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl)
      , (nnet_softmax_layer6_t_result_t_softmax_config7_for_3_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_1_nl)}),
      ({6'b000000 , CALC_SOFTMAX_LOOP_6_or_cse}), {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_644_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_273_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_305_nl)
      , (and_193_nl) , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_652_nl)
      , (and_174_nl) , and_dcpl_175});
  assign and_2658_cse = IndexLoop_stage_0 & IndexLoop_asn_3_itm_1;
  assign nor_668_cse = ~((fsm_output[2:1]!=2'b00));
  assign and_203_m1c = or_dcpl_448 & IndexLoop_stage_0_2;
  assign or_888_cse = (fsm_output[5:4]!=2'b00);
  assign or_647_cse_1 = (fsm_output[3:2]!=2'b00);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_641_cse
      = and_dcpl_207 & and_dcpl_204 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_272_rgt
      = (and_dcpl_200 & and_dcpl_197 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_641_cse;
  assign MultLoop_and_251_rgt = (~ or_dcpl_571) & and_203_m1c & and_dcpl_65;
  assign MultLoop_and_252_rgt = or_dcpl_571 & and_203_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_640_cse
      = and_dcpl_210 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_639_cse
      = (~ IndexLoop_stage_0_2) & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_243_rgt
      = nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_639_cse
      | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_640_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_642_rgt
      = or_dcpl_501 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
      = IndexLoop_stage_0 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_63_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_491_itm)) & (~ nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_243_rgt);
  assign and_215_m1c = or_dcpl_446 & IndexLoop_stage_0_2;
  assign mux_509_cse = MUX_s_1_2_2(mux_tmp_81, or_tmp_48, fsm_output[3]);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_636_cse
      = and_dcpl_219 & and_dcpl_216 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_271_rgt
      = (and_dcpl_212 & and_dcpl_197 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_636_cse;
  assign MultLoop_and_243_rgt = (~ or_dcpl_573) & and_215_m1c & and_dcpl_65;
  assign MultLoop_and_244_rgt = or_dcpl_573 & and_215_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_637_rgt
      = or_dcpl_505 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_64_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_501_itm)) & (~ nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_243_rgt);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_482_m1c
      = nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
      | (~ mux_501_itm);
  assign and_226_m1c = or_dcpl_444 & IndexLoop_stage_0_2;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_65_cse
      = core_wen & (and_dcpl_65 | and_dcpl_60);
  assign and_225_rgt = and_dcpl_200 & and_dcpl_223 & (~ and_dcpl_60);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_304_rgt
      = ((~ or_dcpl_575) & and_226_m1c & (~ and_dcpl_60)) | (and_dcpl_229 & and_dcpl_227
      & and_dcpl_60);
  assign MultLoop_and_242_rgt = or_dcpl_575 & and_226_m1c & (~ and_dcpl_60);
  assign and_232_rgt = or_dcpl_513 & IndexLoop_stage_0_2 & and_dcpl_60;
  assign and_238_m1c = or_dcpl_443 & IndexLoop_stage_0_2;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_629_cse
      = and_dcpl_239 & and_dcpl_204 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_270_rgt
      = (and_dcpl_181 & and_dcpl_235 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_629_cse;
  assign MultLoop_and_239_rgt = (~ or_dcpl_576) & and_238_m1c & and_dcpl_65;
  assign MultLoop_and_240_rgt = or_dcpl_576 & and_238_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_630_rgt
      = or_dcpl_516 & and_dcpl_176 & and_dcpl_60;
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_6_and_seb = reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_1_ftd
      & (~((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_2_reg[4:3]==2'b11)));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_6_nor_2_nl = ~(MUX_v_3_2_2((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_2_reg[2:0]),
      3'b111, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_6_sva_mx0w0));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_6_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl
      = ~(MUX_v_3_2_2((nnet_softmax_layer6_t_result_t_softmax_config7_for_6_nor_2_nl),
      3'b111, nnet_softmax_layer6_t_result_t_softmax_config7_for_6_and_seb));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_6_nor_3_nl = ~(MUX_v_12_2_2(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_3_reg,
      12'b111111111111, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_6_sva_mx0w0));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_6_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_1_nl
      = ~(MUX_v_12_2_2((nnet_softmax_layer6_t_result_t_softmax_config7_for_6_nor_3_nl),
      12'b111111111111, nnet_softmax_layer6_t_result_t_softmax_config7_for_6_and_seb));
  assign and_615_nl = and_dcpl_588 & and_dcpl_573;
  assign and_616_nl = and_dcpl_590 & and_dcpl_573;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_796_rgt
      = MUX1HOT_v_17_7_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_sva_1[16:0]),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_20_sva_1[16:0]),
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0}),
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0}),
      ({2'b00 , (nnet_softmax_layer6_t_result_t_softmax_config7_for_6_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl)
      , (nnet_softmax_layer6_t_result_t_softmax_config7_for_6_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_1_nl)}),
      {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_270_rgt ,
      MultLoop_and_239_rgt , MultLoop_and_240_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_630_rgt
      , (and_615_nl) , (and_616_nl) , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_sva_2_mx0c3});
  assign nor_662_cse = ~((fsm_output[7]) | (~ (fsm_output[0])) | (~ (fsm_output[1]))
      | (fsm_output[2]) | (~ (fsm_output[3])));
  assign or_1875_cse = (fsm_output[1:0]!=2'b00);
  assign and_2657_cse = or_1875_cse & (fsm_output[2]);
  assign and_244_m1c = or_dcpl_442 & IndexLoop_stage_0_2;
  assign and_243_rgt = and_dcpl_212 & and_dcpl_223 & (~ and_dcpl_60);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_303_rgt
      = ((~ or_dcpl_577) & and_244_m1c & (~ and_dcpl_60)) | (and_dcpl_229 & and_dcpl_188
      & and_dcpl_60);
  assign MultLoop_and_238_rgt = or_dcpl_577 & and_244_m1c & (~ and_dcpl_60);
  assign and_246_rgt = or_dcpl_517 & IndexLoop_stage_0_2 & and_dcpl_60;
  assign and_250_m1c = or_dcpl_441 & IndexLoop_stage_0_2;
  assign or_941_cse = (fsm_output[4:3]!=2'b00);
  assign nor_298_cse = ~((fsm_output[4:3]!=2'b00));
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_269_rgt
      = (and_dcpl_247 & and_dcpl_235 & and_dcpl_65) | (and_dcpl_251 & and_dcpl_204
      & and_dcpl_60);
  assign MultLoop_and_235_rgt = (~ or_dcpl_578) & and_250_m1c & and_dcpl_65;
  assign MultLoop_and_236_rgt = or_dcpl_578 & and_250_m1c & and_dcpl_65;
  assign and_254_rgt = or_dcpl_513 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_68_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_533_itm)) & (~ nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_243_rgt);
  assign and_258_m1c = or_dcpl_440 & IndexLoop_stage_0_2;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_268_rgt
      = (and_dcpl_255 & and_dcpl_197 & (~ and_dcpl_60)) | (and_dcpl_218 & (~ (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[4]))
      & and_dcpl_227 & and_dcpl_60);
  assign MultLoop_and_233_rgt = (~ or_dcpl_579) & and_258_m1c & (~ and_dcpl_60);
  assign MultLoop_and_234_rgt = or_dcpl_579 & and_258_m1c & (~ and_dcpl_60);
  assign and_261_rgt = or_dcpl_518 & IndexLoop_stage_0_2 & and_dcpl_60;
  assign and_266_m1c = or_dcpl_439 & IndexLoop_stage_0_2;
  assign and_265_rgt = and_dcpl_263 & and_dcpl_261 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_302_rgt
      = ((~ or_dcpl_580) & and_266_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_641_cse;
  assign MultLoop_and_232_rgt = or_dcpl_580 & and_266_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_70_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_544_itm)) & (~ nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_243_rgt);
  assign and_269_m1c = or_dcpl_438 & IndexLoop_stage_0_2;
  assign and_268_rgt = and_dcpl_266 & and_dcpl_197 & (~ and_dcpl_60);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_301_rgt
      = ((~ or_dcpl_581) & and_269_m1c & (~ and_dcpl_60)) | (and_dcpl_206 & (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[4])
      & (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[1])
      & (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[0])
      & IndexLoop_stage_0_2 & and_dcpl_60);
  assign MultLoop_and_230_rgt = or_dcpl_581 & and_269_m1c & (~ and_dcpl_60);
  assign and_274_rgt = or_dcpl_520 & IndexLoop_stage_0_2 & and_dcpl_60;
  assign and_277_m1c = or_dcpl_437 & IndexLoop_stage_0_2;
  assign mux_389_cse = MUX_s_1_2_2(or_611_cse, mux_tmp_377, fsm_output[2]);
  assign and_276_rgt = and_dcpl_274 & and_dcpl_261 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_300_rgt
      = ((~ or_dcpl_582) & and_277_m1c & and_dcpl_65) | (and_dcpl_277 & and_dcpl_204
      & and_dcpl_60);
  assign MultLoop_and_228_rgt = or_dcpl_582 & and_277_m1c & and_dcpl_65;
  assign and_280_rgt = or_dcpl_522 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_72_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_556_itm)) & (~ nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_243_rgt);
  assign and_283_m1c = or_dcpl_436 & IndexLoop_stage_0_2;
  assign mux_425_cse = MUX_s_1_2_2(nand_tmp_14, or_1298_cse, fsm_output[1]);
  assign and_282_rgt = and_dcpl_255 & and_dcpl_223 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_607_cse
      = and_dcpl_283 & and_dcpl_204 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_299_rgt
      = ((~ or_dcpl_583) & and_283_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_607_cse;
  assign MultLoop_and_226_rgt = or_dcpl_583 & and_283_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_608_rgt
      = or_dcpl_525 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_73_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_sva_2_mx0c2)
      & (~ nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_243_rgt);
  assign and_288_m1c = or_dcpl_435 & IndexLoop_stage_0_2;
  assign and_287_rgt = and_dcpl_263 & and_dcpl_235 & (~ and_dcpl_60);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_298_rgt
      = ((~ or_dcpl_584) & and_288_m1c & (~ and_dcpl_60)) | (and_dcpl_229 & (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[1:0]==2'b00)
      & IndexLoop_stage_0_2 & and_dcpl_60);
  assign MultLoop_and_224_rgt = or_dcpl_584 & and_288_m1c & (~ and_dcpl_60);
  assign and_292_rgt = or_dcpl_526 & IndexLoop_stage_0_2 & and_dcpl_60;
  assign and_295_m1c = or_dcpl_434 & IndexLoop_stage_0_2;
  assign and_294_rgt = and_dcpl_266 & and_dcpl_223 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_600_cse
      = and_dcpl_295 & and_dcpl_216 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_297_rgt
      = ((~ or_dcpl_585) & and_295_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_600_cse;
  assign MultLoop_and_222_rgt = or_dcpl_585 & and_295_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_601_rgt
      = or_dcpl_528 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_75_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_sva_2_mx0c2)
      & (~ nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_243_rgt);
  assign and_300_m1c = or_dcpl_433 & IndexLoop_stage_0_2;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_595_cse
      = and_dcpl_207 & and_dcpl_216 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_267_rgt
      = (and_dcpl_274 & and_dcpl_235 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_595_cse;
  assign MultLoop_and_219_rgt = (~ or_dcpl_586) & and_300_m1c & and_dcpl_65;
  assign MultLoop_and_220_rgt = or_dcpl_586 & and_300_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_596_rgt
      = or_dcpl_529 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_76_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_571_itm)) & (~ nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_243_rgt);
  assign and_306_m1c = or_dcpl_432 & IndexLoop_stage_0_2;
  assign and_305_rgt = and_dcpl_303 & and_dcpl_197 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_591_cse
      = and_dcpl_295 & and_dcpl_204 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_296_rgt
      = ((~ or_dcpl_587) & and_306_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_591_cse;
  assign MultLoop_and_218_rgt = or_dcpl_587 & and_306_m1c & and_dcpl_65;
  assign and_308_rgt = or_dcpl_531 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_77_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_sva_2_mx0c2)
      & (~ nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_243_rgt);
  assign and_312_m1c = or_dcpl_430 & IndexLoop_stage_0_2;
  assign and_311_rgt = and_dcpl_309 & and_dcpl_197 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_586_cse
      = and_dcpl_312 & and_dcpl_216 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_295_rgt
      = ((~ or_dcpl_589) & and_312_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_586_cse;
  assign MultLoop_and_214_rgt = or_dcpl_589 & and_312_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_587_rgt
      = or_dcpl_533 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_78_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_sva_2_mx0c2)
      & (~ nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_243_rgt);
  assign and_317_m1c = or_dcpl_428 & IndexLoop_stage_0_2;
  assign or_1405_cse = (fsm_output[5:3]!=3'b000);
  assign and_316_rgt = and_dcpl_303 & and_dcpl_223 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_581_cse
      = and_dcpl_312 & and_dcpl_204 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_294_rgt
      = ((~ or_dcpl_591) & and_317_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_581_cse;
  assign MultLoop_and_210_rgt = or_dcpl_591 & and_317_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_582_rgt
      = or_dcpl_534 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_79_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_588_itm)) & (~ nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_243_rgt);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_472_m1c
      = nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
      | (~ mux_588_itm);
  assign and_321_m1c = or_dcpl_426 & IndexLoop_stage_0_2;
  assign and_320_rgt = and_dcpl_309 & and_dcpl_223 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_576_cse
      = and_dcpl_239 & and_dcpl_216 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_293_rgt
      = ((~ or_dcpl_593) & and_321_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_576_cse;
  assign MultLoop_and_208_rgt = or_dcpl_593 & and_321_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_577_rgt
      = or_dcpl_535 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_80_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_595_itm)) & (~ nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_243_rgt);
  assign and_329_m1c = or_dcpl_425 & and_dcpl_176;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_conc_231_itm_11_0
      = MUX_v_12_2_2(CALC_SOFTMAX_LOOP_6_or_cse, ({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_4_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd_2}),
      and_dcpl_338);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_570_cse
      = and_dcpl_329 & and_dcpl_204 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_266_rgt
      = (and_dcpl_326 & and_dcpl_325 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_570_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_307_rgt
      = ((~ or_dcpl_594) & and_329_m1c & and_dcpl_65) | (and_dcpl_176 & MultLoop_2_and_5_itm_1
      & and_dcpl_55);
  assign MultLoop_and_206_rgt = or_dcpl_594 & and_329_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_566_rgt
      = IndexLoop_stage_0 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_569_cse
      = and_dcpl_210 & and_dcpl_55;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_567_cse
      = and_dcpl_210 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_571_rgt
      = or_dcpl_537 & and_dcpl_176 & and_dcpl_60;
  assign and_334_rgt = and_dcpl_176 & (~ MultLoop_2_and_5_itm_1) & and_dcpl_55;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_946_rgt
      = and_dcpl_588 & and_dcpl_154;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_948_rgt
      = and_dcpl_590 & and_dcpl_154;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_745_rgt
      = MUX1HOT_v_7_8_2((z_out_20[16:10]), (z_out_21[16:10]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_sva_1[16:10]),
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12
      , (nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0[11:10])}),
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_10}),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_12_sva_1[16:10]),
      (nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_3_sva_1[16:10]),
      ({5'b00000 , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_conc_231_itm_11_0[11:10])}),
      {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_266_rgt ,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_307_rgt , MultLoop_and_206_rgt
      , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_946_rgt
      , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_948_rgt
      , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_571_rgt
      , and_334_rgt , and_dcpl_324});
  assign and_2654_cse = (z_out_23_22_8[10]) & (fsm_output[6]);
  assign nor_654_cse = ~((~ (fsm_output[4])) | (~ (fsm_output[7])) | (fsm_output[6])
      | (fsm_output[2]) | (~ (fsm_output[1])) | (fsm_output[0]));
  assign nand_209_cse = ~((fsm_output[1:0]==2'b11));
  assign nand_210_cse = ~((fsm_output[2:0]==3'b111));
  assign nor_649_cse = ~((fsm_output[2]) | nand_209_cse);
  assign or_1876_cse = (~ or_tmp_940) | (fsm_output[4]);
  assign and_337_m1c = or_dcpl_424 & IndexLoop_stage_0_2;
  assign and_336_rgt = and_dcpl_334 & and_dcpl_197 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_292_rgt
      = ((~ or_dcpl_595) & and_337_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_629_cse;
  assign MultLoop_and_204_rgt = or_dcpl_595 & and_337_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse
      = ~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_639_cse
      | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_640_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_82_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_616_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_342_m1c = or_dcpl_423 & IndexLoop_stage_0_2;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_557_cse
      = and_dcpl_329 & and_dcpl_216 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_265_rgt
      = (and_dcpl_339 & and_dcpl_261 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_557_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_306_rgt
      = ((~ or_dcpl_596) & and_342_m1c & and_dcpl_65) | (and_dcpl_194 & (ReuseLoop_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_outidx_const_assign_1_ReuseLoop_2_asn_tmp_3_2_0_psp_sva_1[2:1]==2'b10)
      & and_dcpl_55);
  assign MultLoop_and_202_rgt = or_dcpl_596 & and_342_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_558_rgt
      = or_dcpl_538 & and_dcpl_176 & and_dcpl_60;
  assign and_347_rgt = or_dcpl_540 & and_dcpl_176 & and_dcpl_55;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_136_cse
      = ~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_639_cse
      | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_640_cse
      | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_569_cse);
  assign and_599_nl = and_dcpl_588 & and_dcpl_62;
  assign and_600_nl = and_dcpl_590 & and_dcpl_62;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_747_rgt
      = MUX1HOT_v_17_8_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_sva_1[16:0]),
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0}),
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0}),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_13_sva_1[16:0]),
      (nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_4_sva_1[16:0]),
      ({5'b00000 , CALC_SOFTMAX_LOOP_6_or_cse}), {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_265_rgt
      , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_306_rgt ,
      MultLoop_and_202_rgt , (and_599_nl) , (and_600_nl) , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_558_rgt
      , and_347_rgt , and_dcpl_338});
  assign and_350_m1c = or_dcpl_422 & IndexLoop_stage_0_2;
  assign and_349_rgt = and_dcpl_347 & and_dcpl_197 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_551_cse
      = and_dcpl_277 & and_dcpl_216 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_291_rgt
      = ((~ or_dcpl_597) & and_350_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_551_cse;
  assign MultLoop_and_200_rgt = or_dcpl_597 & and_350_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_552_rgt
      = or_dcpl_541 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_84_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_631_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_357_m1c = or_dcpl_421 & IndexLoop_stage_0_2;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_545_cse
      = and_dcpl_357 & and_dcpl_204 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_264_rgt
      = (and_dcpl_354 & and_dcpl_261 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_545_cse
      | (and_dcpl_194 & (~ (ReuseLoop_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_outidx_const_assign_1_ReuseLoop_2_asn_tmp_3_2_0_psp_sva_1[1]))
      & nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_out_index_3_0_sva_1_2
      & and_dcpl_55);
  assign MultLoop_and_197_rgt = (~ or_dcpl_598) & and_357_m1c & and_dcpl_65;
  assign MultLoop_and_198_rgt = or_dcpl_598 & and_357_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_546_rgt
      = or_dcpl_543 & and_dcpl_176 & and_dcpl_60;
  assign and_363_rgt = or_dcpl_544 & and_dcpl_176 & and_dcpl_55;
  assign and_601_nl = and_dcpl_588 & and_dcpl_157;
  assign and_602_nl = and_dcpl_590 & and_dcpl_157;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_748_rgt
      = MUX1HOT_v_17_8_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_sva_1[16:0]),
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0}),
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0}),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_14_sva_1[16:0]),
      (nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_5_sva_1[16:0]),
      ({5'b00000 , CALC_SOFTMAX_LOOP_6_or_cse}), {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_264_rgt
      , MultLoop_and_197_rgt , MultLoop_and_198_rgt , (and_601_nl) , (and_602_nl)
      , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_546_rgt
      , and_363_rgt , and_dcpl_353});
  assign or_1637_cse = (~ (fsm_output[0])) | (~ IndexLoop_stage_0_2) | (fsm_output[3:2]!=2'b00);
  assign nor_642_cse = ~((fsm_output[7]) | (~ (fsm_output[0])) | (~ IndexLoop_stage_0_2)
      | IndexLoop_stage_0 | (fsm_output[3:2]!=2'b01));
  assign nor_647_cse = ~((fsm_output[6]) | (fsm_output[4]) | (~ (fsm_output[0]))
      | (~ IndexLoop_stage_0_2) | IndexLoop_stage_0 | (~ (fsm_output[2])));
  assign nor_646_cse = ~((fsm_output[6]) | (fsm_output[4]) | (~ (fsm_output[0]))
      | (~ IndexLoop_stage_0_2) | (fsm_output[2]));
  assign and_365_m1c = or_dcpl_420 & IndexLoop_stage_0_2;
  assign or_611_cse = (fsm_output[5:3]!=3'b000) | mux_661_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_539_cse
      = and_dcpl_365 & and_dcpl_216 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_263_rgt
      = (and_dcpl_334 & and_dcpl_223 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_539_cse;
  assign MultLoop_and_195_rgt = (~ or_dcpl_599) & and_365_m1c & and_dcpl_65;
  assign MultLoop_and_196_rgt = or_dcpl_599 & and_365_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_540_rgt
      = or_dcpl_545 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_86_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_643_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_372_m1c = or_dcpl_419 & IndexLoop_stage_0_2;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_533_cse
      = and_dcpl_357 & and_dcpl_216 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_262_rgt
      = (and_dcpl_339 & and_dcpl_235 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_533_cse
      | (and_dcpl_176 & MultLoop_2_and_14_itm_1 & and_dcpl_55);
  assign MultLoop_and_193_rgt = (~ or_dcpl_600) & and_372_m1c & and_dcpl_65;
  assign MultLoop_and_194_rgt = or_dcpl_600 & and_372_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_534_rgt
      = or_dcpl_546 & and_dcpl_176 & and_dcpl_60;
  assign and_376_rgt = and_dcpl_176 & (~ MultLoop_2_and_14_itm_1) & and_dcpl_55;
  assign and_603_nl = and_dcpl_588 & and_dcpl_57;
  assign and_604_nl = and_dcpl_590 & and_dcpl_57;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_749_rgt
      = MUX1HOT_v_17_8_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_sva_1[16:0]),
      nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0}),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_15_sva_1[16:0]),
      (nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_6_sva_1[16:0]),
      ({5'b00000 , CALC_SOFTMAX_LOOP_6_or_cse}), {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_262_rgt
      , MultLoop_and_193_rgt , MultLoop_and_194_rgt , (and_603_nl) , (and_604_nl)
      , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_534_rgt
      , and_376_rgt , and_dcpl_369});
  assign and_2650_cse = (fsm_output[3:2]==2'b11);
  assign and_378_m1c = or_dcpl_418 & IndexLoop_stage_0_2;
  assign and_377_rgt = and_dcpl_347 & and_dcpl_223 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_527_cse
      = and_dcpl_378 & and_dcpl_216 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_290_rgt
      = ((~ or_dcpl_601) & and_378_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_527_cse;
  assign MultLoop_and_192_rgt = or_dcpl_601 & and_378_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_528_rgt
      = or_dcpl_547 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_88_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_654_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_383_m1c = or_dcpl_417 & IndexLoop_stage_0_2;
  assign mux_661_cse = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), fsm_output[6]);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_521_cse
      = and_dcpl_378 & and_dcpl_204 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_261_rgt
      = (and_dcpl_354 & and_dcpl_235 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_521_cse
      | (and_dcpl_176 & MultLoop_2_and_15_itm_1 & and_dcpl_55);
  assign MultLoop_and_189_rgt = (~ or_dcpl_602) & and_383_m1c & and_dcpl_65;
  assign MultLoop_and_190_rgt = or_dcpl_602 & and_383_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_522_rgt
      = or_dcpl_548 & and_dcpl_176 & and_dcpl_60;
  assign and_387_rgt = and_dcpl_176 & (~ MultLoop_2_and_15_itm_1) & and_dcpl_55;
  assign nor_959_cse = ~((fsm_output[3]) | (fsm_output[5]));
  assign and_389_m1c = or_dcpl_416 & IndexLoop_stage_0_2;
  assign and_388_rgt = and_dcpl_354 & and_dcpl_197 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_289_rgt
      = ((~ or_dcpl_602) & and_389_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_521_cse;
  assign MultLoop_and_188_rgt = or_dcpl_602 & and_389_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_90_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_665_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_391_m1c = or_dcpl_415 & IndexLoop_stage_0_2;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_260_rgt
      = (and_dcpl_347 & and_dcpl_261 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_527_cse
      | (and_dcpl_176 & MultLoop_2_MultLoop_2_nor_2_itm_1 & and_dcpl_55);
  assign MultLoop_and_185_rgt = (~ or_dcpl_601) & and_391_m1c & and_dcpl_65;
  assign MultLoop_and_186_rgt = or_dcpl_601 & and_391_m1c & and_dcpl_65;
  assign and_393_rgt = and_dcpl_176 & (~ MultLoop_2_MultLoop_2_nor_2_itm_1) & and_dcpl_55;
  assign and_395_m1c = or_dcpl_414 & IndexLoop_stage_0_2;
  assign and_394_rgt = and_dcpl_339 & and_dcpl_197 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_288_rgt
      = ((~ or_dcpl_600) & and_395_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_533_cse;
  assign MultLoop_and_184_rgt = or_dcpl_600 & and_395_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_92_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_681_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_397_m1c = or_dcpl_413 & IndexLoop_stage_0_2;
  assign or_1419_tmp = or_dcpl_539 | nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_out_index_3_0_sva_1_2;
  assign or_1083_nl = nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_out_index_3_0_sva_1_2
      | (ReuseLoop_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_outidx_const_assign_1_ReuseLoop_2_asn_tmp_3_2_0_psp_sva_1[1:0]!=2'b00);
  assign mux_690_nl = MUX_s_1_2_2(and_2658_cse, or_tmp_384, or_1083_nl);
  assign or_1084_tmp = (or_1419_tmp & and_dcpl_185) | (mux_690_nl) | (~ IndexLoop_stage_0_2);
  assign and_404_m1c = or_dcpl_412 & IndexLoop_stage_0_2;
  assign and_403_rgt = and_dcpl_354 & and_dcpl_223 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_287_rgt
      = ((~ or_dcpl_598) & and_404_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_545_cse;
  assign MultLoop_and_180_rgt = or_dcpl_598 & and_404_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_94_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_692_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_408_m1c = or_dcpl_411 & IndexLoop_stage_0_2;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_258_rgt
      = (and_dcpl_347 & and_dcpl_235 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_551_cse;
  assign MultLoop_and_177_rgt = (~ or_dcpl_597) & and_408_m1c & and_dcpl_65;
  assign MultLoop_and_178_rgt = or_dcpl_597 & and_408_m1c & and_dcpl_65;
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_4_and_seb = reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd
      & (~((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_2_reg[4:3]==2'b11)));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_4_nor_2_nl = ~(MUX_v_3_2_2((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_2_reg[2:0]),
      3'b111, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_4_sva_mx0w1));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_4_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl
      = ~(MUX_v_3_2_2((nnet_softmax_layer6_t_result_t_softmax_config7_for_4_nor_2_nl),
      3'b111, nnet_softmax_layer6_t_result_t_softmax_config7_for_4_and_seb));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_4_nor_3_nl = ~(MUX_v_2_2_2(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_4_reg,
      2'b11, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_4_sva_mx0w1));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_4_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_1_nl
      = ~(MUX_v_2_2_2((nnet_softmax_layer6_t_result_t_softmax_config7_for_4_nor_3_nl),
      2'b11, nnet_softmax_layer6_t_result_t_softmax_config7_for_4_and_seb));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_4_nor_4_nl = ~(MUX_v_10_2_2(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd_2,
      10'b1111111111, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_4_sva_mx0w1));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_4_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_2_nl
      = ~(MUX_v_10_2_2((nnet_softmax_layer6_t_result_t_softmax_config7_for_4_nor_4_nl),
      10'b1111111111, nnet_softmax_layer6_t_result_t_softmax_config7_for_4_and_seb));
  assign and_611_nl = and_dcpl_588 & and_dcpl_567;
  assign and_612_nl = and_dcpl_590 & and_dcpl_567;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_778_rgt
      = MUX1HOT_v_17_7_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_sva_1[16:0]),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_19_sva_1[16:0]),
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_16_0_lpi_1_dfm_mx0w2_16_15
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_16_0_lpi_1_dfm_mx0w2_14_0}),
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0}),
      ({2'b00 , (nnet_softmax_layer6_t_result_t_softmax_config7_for_4_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl)
      , (nnet_softmax_layer6_t_result_t_softmax_config7_for_4_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_1_nl)
      , (nnet_softmax_layer6_t_result_t_softmax_config7_for_4_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_2_nl)}),
      {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_258_rgt ,
      MultLoop_and_177_rgt , MultLoop_and_178_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_552_rgt
      , (and_611_nl) , (and_612_nl) , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_sva_2_mx0c3});
  assign nor_622_cse = ~((fsm_output[0]) | (fsm_output[4]) | (fsm_output[6]) | (~
      (fsm_output[3])) | (fsm_output[2]) | (fsm_output[1]));
  assign and_410_m1c = or_dcpl_410 & IndexLoop_stage_0_2;
  assign and_409_rgt = and_dcpl_339 & and_dcpl_223 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_286_rgt
      = ((~ or_dcpl_596) & and_410_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_557_cse;
  assign MultLoop_and_176_rgt = or_dcpl_596 & and_410_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_96_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_703_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_415_m1c = or_dcpl_409 & IndexLoop_stage_0_2;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_479_cse
      = and_dcpl_415 & and_dcpl_204 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_257_rgt
      = (and_dcpl_334 & and_dcpl_235 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_479_cse;
  assign MultLoop_and_173_rgt = (~ or_dcpl_595) & and_415_m1c & and_dcpl_65;
  assign MultLoop_and_174_rgt = or_dcpl_595 & and_415_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_480_rgt
      = or_dcpl_551 & and_dcpl_176 & and_dcpl_60;
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_5_and_seb = reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_1_ftd
      & (~((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_2_reg[4:3]==2'b11)));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_5_nor_2_nl = ~(MUX_v_3_2_2((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_2_reg[2:0]),
      3'b111, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_5_sva_mx0w0));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_5_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl
      = ~(MUX_v_3_2_2((nnet_softmax_layer6_t_result_t_softmax_config7_for_5_nor_2_nl),
      3'b111, nnet_softmax_layer6_t_result_t_softmax_config7_for_5_and_seb));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_5_nor_3_nl = ~(MUX_v_12_2_2(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_3_reg,
      12'b111111111111, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_5_sva_mx0w0));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_5_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_1_nl
      = ~(MUX_v_12_2_2((nnet_softmax_layer6_t_result_t_softmax_config7_for_5_nor_3_nl),
      12'b111111111111, nnet_softmax_layer6_t_result_t_softmax_config7_for_5_and_seb));
  assign and_613_nl = and_dcpl_588 & and_dcpl_570;
  assign and_614_nl = and_dcpl_590 & and_dcpl_570;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_776_rgt
      = MUX1HOT_v_17_7_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_sva_1[16:0]),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_2_sva_1[16:0]),
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0}),
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0}),
      ({2'b00 , (nnet_softmax_layer6_t_result_t_softmax_config7_for_5_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl)
      , (nnet_softmax_layer6_t_result_t_softmax_config7_for_5_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_1_nl)}),
      {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_257_rgt ,
      MultLoop_and_173_rgt , MultLoop_and_174_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_480_rgt
      , (and_613_nl) , (and_614_nl) , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_sva_2_mx0c3});
  assign and_420_m1c = or_dcpl_408 & IndexLoop_stage_0_2;
  assign and_419_rgt = and_dcpl_326 & and_dcpl_197 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_285_rgt
      = ((~ or_dcpl_594) & and_420_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_570_cse;
  assign MultLoop_and_172_rgt = or_dcpl_594 & and_420_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_98_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_714_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_424_m1c = or_dcpl_407 & IndexLoop_stage_0_2;
  assign nand_52_cse = ~((fsm_output[2:1]==2'b11));
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_256_rgt
      = (and_dcpl_309 & and_dcpl_261 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_576_cse;
  assign MultLoop_and_169_rgt = (~ or_dcpl_593) & and_424_m1c & and_dcpl_65;
  assign MultLoop_and_170_rgt = or_dcpl_593 & and_424_m1c & and_dcpl_65;
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_7_and_seb = reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_1_ftd
      & (~((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_2_reg[4:3]==2'b11)));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_7_nor_2_nl = ~(MUX_v_3_2_2((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_2_reg[2:0]),
      3'b111, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_7_sva_mx0w0));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_7_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl
      = ~(MUX_v_3_2_2((nnet_softmax_layer6_t_result_t_softmax_config7_for_7_nor_2_nl),
      3'b111, nnet_softmax_layer6_t_result_t_softmax_config7_for_7_and_seb));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_7_nor_3_nl = ~(MUX_v_12_2_2(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_3_reg,
      12'b111111111111, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_7_sva_mx0w0));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_7_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_1_nl
      = ~(MUX_v_12_2_2((nnet_softmax_layer6_t_result_t_softmax_config7_for_7_nor_3_nl),
      12'b111111111111, nnet_softmax_layer6_t_result_t_softmax_config7_for_7_and_seb));
  assign and_617_nl = and_dcpl_588 & and_dcpl_576;
  assign and_618_nl = and_dcpl_590 & and_dcpl_576;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_774_rgt
      = MUX1HOT_v_17_7_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_sva_1[16:0]),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_21_sva_1[16:0]),
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0}),
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0}),
      ({2'b00 , (nnet_softmax_layer6_t_result_t_softmax_config7_for_7_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl)
      , (nnet_softmax_layer6_t_result_t_softmax_config7_for_7_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_1_nl)}),
      {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_256_rgt ,
      MultLoop_and_169_rgt , MultLoop_and_170_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_577_rgt
      , (and_617_nl) , (and_618_nl) , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_sva_2_mx0c3});
  assign nor_610_cse = ~((fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[7])
      | (fsm_output[0]) | (~ (fsm_output[3])));
  assign and_427_m1c = or_dcpl_406 & IndexLoop_stage_0_2;
  assign and_426_rgt = and_dcpl_424 & and_dcpl_197 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_465_cse
      = and_dcpl_427 & and_dcpl_216 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_284_rgt
      = ((~ or_dcpl_592) & and_427_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_465_cse;
  assign MultLoop_and_168_rgt = or_dcpl_592 & and_427_m1c & and_dcpl_65;
  assign and_430_rgt = or_dcpl_552 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_100_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_725_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_434_m1c = or_dcpl_405 & IndexLoop_stage_0_2;
  assign and_862_cse = (fsm_output[4:3]==2'b11);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_255_rgt
      = (and_dcpl_303 & and_dcpl_261 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_581_cse;
  assign MultLoop_and_165_rgt = (~ or_dcpl_591) & and_434_m1c & and_dcpl_65;
  assign MultLoop_and_166_rgt = or_dcpl_591 & and_434_m1c & and_dcpl_65;
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_8_nor_2_nl = ~(MUX_v_15_2_2((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd_1[14:0]),
      15'b111111111111111, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_8_sva_mx0w0));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_8_and_nl = reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd
      & (~((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd_1[16:15]==2'b11)));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_8_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl
      = ~(MUX_v_15_2_2((nnet_softmax_layer6_t_result_t_softmax_config7_for_8_nor_2_nl),
      15'b111111111111111, (nnet_softmax_layer6_t_result_t_softmax_config7_for_8_and_nl)));
  assign and_619_nl = and_dcpl_588 & and_dcpl_579;
  assign and_620_nl = and_dcpl_590 & and_dcpl_579;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_772_rgt
      = MUX1HOT_v_17_7_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_sva_1[16:0]),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_22_sva_1[16:0]),
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_12
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0}),
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0}),
      ({2'b00 , (nnet_softmax_layer6_t_result_t_softmax_config7_for_8_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl)}),
      {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_255_rgt ,
      MultLoop_and_165_rgt , MultLoop_and_166_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_582_rgt
      , (and_619_nl) , (and_620_nl) , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_sva_2_mx0c3});
  assign and_2642_cse = (fsm_output[2:0]==3'b111);
  assign nor_601_nl = ~((fsm_output[4]) | (fsm_output[2]) | nand_209_cse);
  assign nor_602_nl = ~(IndexLoop_stage_0 | (fsm_output[4]) | (~ (fsm_output[2]))
      | (~ (fsm_output[0])) | (fsm_output[1]));
  assign mux_1161_nl = MUX_s_1_2_2((nor_601_nl), (nor_602_nl), fsm_output[6]);
  assign and_2640_nl = IndexLoop_stage_0_2 & (mux_1161_nl);
  assign and_2641_nl = (fsm_output[4]) & (fsm_output[2]) & (fsm_output[0]) & (~ (fsm_output[1]));
  assign mux_1162_cse = MUX_s_1_2_2((and_2640_nl), (and_2641_nl), fsm_output[3]);
  assign and_436_m1c = or_dcpl_404 & IndexLoop_stage_0_2;
  assign and_435_rgt = and_dcpl_326 & and_dcpl_223 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_456_cse
      = and_dcpl_427 & and_dcpl_204 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_283_rgt
      = ((~ or_dcpl_590) & and_436_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_456_cse;
  assign MultLoop_and_164_rgt = or_dcpl_590 & and_436_m1c & and_dcpl_65;
  assign and_438_rgt = or_dcpl_554 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_102_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_739_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_441_m1c = or_dcpl_402 & IndexLoop_stage_0_2;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_254_rgt
      = (and_dcpl_309 & and_dcpl_235 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_586_cse;
  assign MultLoop_and_161_rgt = (~ or_dcpl_589) & and_441_m1c & and_dcpl_65;
  assign MultLoop_and_162_rgt = or_dcpl_589 & and_441_m1c & and_dcpl_65;
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_9_nor_2_nl = ~(MUX_v_15_2_2((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd_1[14:0]),
      15'b111111111111111, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_9_sva_mx0w0));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_9_and_nl = reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd
      & (~((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd_1[16:15]==2'b11)));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_9_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl
      = ~(MUX_v_15_2_2((nnet_softmax_layer6_t_result_t_softmax_config7_for_9_nor_2_nl),
      15'b111111111111111, (nnet_softmax_layer6_t_result_t_softmax_config7_for_9_and_nl)));
  assign and_621_nl = and_dcpl_588 & and_dcpl_517;
  assign and_622_nl = and_dcpl_590 & and_dcpl_517;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_770_rgt
      = MUX1HOT_v_17_7_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_sva_1[16:0]),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_23_sva_1[16:0]),
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_12
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_10_0}),
      ({nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_12
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0}),
      ({2'b00 , (nnet_softmax_layer6_t_result_t_softmax_config7_for_9_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl)}),
      {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_254_rgt ,
      MultLoop_and_161_rgt , MultLoop_and_162_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_587_rgt
      , (and_621_nl) , (and_622_nl) , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_sva_2_mx0c3});
  assign and_443_m1c = or_dcpl_400 & IndexLoop_stage_0_2;
  assign and_442_rgt = and_dcpl_424 & and_dcpl_223 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_282_rgt
      = ((~ or_dcpl_588) & and_443_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_595_cse;
  assign MultLoop_and_160_rgt = or_dcpl_588 & and_443_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_104_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_753_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_457_m1c = or_dcpl_398 & and_dcpl_176;
  assign or_10_cse = (fsm_output[2:1]!=2'b00);
  assign or_9_nl = (fsm_output[4]) | (fsm_output[7]);
  assign mux_cse = MUX_s_1_2_2((or_9_nl), or_tmp_2, fsm_output[3]);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_253_rgt
      = (and_dcpl_303 & and_dcpl_325 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_591_cse;
  assign MultLoop_and_157_rgt = (~ or_dcpl_587) & and_457_m1c & and_dcpl_65;
  assign MultLoop_and_158_rgt = or_dcpl_587 & and_457_m1c & and_dcpl_65;
  assign or_1286_cse = (fsm_output[2:1]!=2'b01);
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_10_nor_2_nl = ~(MUX_v_15_2_2((nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2[14:0]),
      15'b111111111111111, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_sva_mx0w0));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_10_and_nl = (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2[17])
      & (~((nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2[16:15]==2'b11)));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_10_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl
      = ~(MUX_v_15_2_2((nnet_softmax_layer6_t_result_t_softmax_config7_for_10_nor_2_nl),
      15'b111111111111111, (nnet_softmax_layer6_t_result_t_softmax_config7_for_10_and_nl)));
  assign IndexLoop_ir_IndexLoop_ir_mux_nl = MUX_v_15_2_2((z_out_13[14:0]), (nnet_softmax_layer6_t_result_t_softmax_config7_for_10_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl),
      and_dcpl_520);
  assign mux_5_nl = MUX_s_1_2_2(mux_tmp_2, or_tmp_1, or_10_cse);
  assign mux_885_nl = MUX_s_1_2_2(mux_cse, or_tmp_1, or_1286_cse);
  assign mux_887_nl = MUX_s_1_2_2((mux_5_nl), (mux_885_nl), fsm_output[0]);
  assign nor_372_nl = ~((mux_887_nl) | or_1398_cse);
  assign IndexLoop_ir_asn_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_3_14_IndexLoop_ir_and_nl
      = MUX_v_15_2_2(15'b000000000000000, (IndexLoop_ir_IndexLoop_ir_mux_nl), (nor_372_nl));
  assign MultLoop_1_1_MultLoop_1_mux_1_nl = MUX_v_15_64_2(({layer3_out_0_16_0_lpi_1_dfm_14_12
      , layer3_out_0_16_0_lpi_1_dfm_11_0}), ({(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_16_0_lpi_1_dfm_16_12[2:0])
      , nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_16_0_lpi_1_dfm_11_0}),
      reg_nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_16_0_lpi_1_dfm_ftd_1,
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_16_0_lpi_1_dfm[14:0]),
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_16_0_lpi_1_dfm[14:0]),
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_16_0_lpi_1_dfm[14:0]),
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_16_0_lpi_1_dfm[14:0]),
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_16_0_lpi_1_dfm[14:0]),
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_16_0_lpi_1_dfm[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_63_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_1_ftd_1[14:0]),
      ({(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_2_reg[2:0])
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_4_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd_2}),
      ({(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_2_reg[2:0])
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_3_reg}),
      ({(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_2_reg[2:0])
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_3_reg}),
      ({(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_2_reg[2:0])
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_3_reg}),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd_1[14:0]),
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_16_0_lpi_1_dfm[14:0]),
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_14_0,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_14_0,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_14_0,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_14_0,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_14_0,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_14_0,
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_16_0_lpi_1_dfm[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_1_ftd_1[14:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_1_ftd_1[14:0]),
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_16_0_lpi_1_dfm[14:0]),
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_16_0_lpi_1_dfm[14:0]),
      InitAccumLoop_1_iacc_6_0_sva_5_0);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_484_nl =
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_2_mx0c0
      | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_566_rgt;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_799_rgt
      = MUX1HOT_v_15_7_2((IndexLoop_ir_asn_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_3_14_IndexLoop_ir_and_nl),
      (z_out_20[14:0]), (z_out_21[14:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_1[14:0]),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_24_sva_1[14:0]),
      (MultLoop_1_1_MultLoop_1_mux_1_nl), ({3'b000 , CALC_SOFTMAX_LOOP_6_or_cse}),
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_484_nl) ,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_253_rgt , MultLoop_and_157_rgt
      , MultLoop_and_158_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_2_mx0c3
      , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_2_mx0c4
      , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_2_mx0c5});
  assign nor_586_cse = ~((fsm_output[7:6]!=2'b10));
  assign and_459_m1c = or_dcpl_396 & IndexLoop_stage_0_2;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_439_cse
      = and_dcpl_365 & and_dcpl_204 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_252_rgt
      = (and_dcpl_274 & and_dcpl_197 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_439_cse;
  assign MultLoop_and_155_rgt = (~ or_dcpl_586) & and_459_m1c & and_dcpl_65;
  assign MultLoop_and_156_rgt = or_dcpl_586 & and_459_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_440_rgt
      = or_dcpl_556 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_106_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_775_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_447_m1c
      = nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
      | (~ mux_775_itm);
  assign and_470_m1c = or_dcpl_395 & and_dcpl_176;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_251_rgt
      = (and_dcpl_266 & and_dcpl_178 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_600_cse;
  assign MultLoop_and_153_rgt = (~ or_dcpl_585) & and_470_m1c & and_dcpl_65;
  assign MultLoop_and_154_rgt = or_dcpl_585 & and_470_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_107_ssc
      = core_wen & (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_2_mx0c0
      | and_dcpl_65 | and_dcpl_158 | and_dcpl_60 | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_2_mx0c4
      | and_dcpl_467) & (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_567_cse
      | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_640_cse));
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_444_cse
      = nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_2_mx0c0
      | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_566_rgt;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_766_rgt
      = MUX1HOT_v_4_6_2((nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_3_14_0[14:11]),
      (z_out_20[14:11]), (z_out_21[14:11]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_1[14:11]),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_25_sva_1[14:11]),
      ({3'b000 , (CALC_SOFTMAX_LOOP_6_or_cse[11])}), {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_444_cse
      , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_251_rgt ,
      MultLoop_and_153_rgt , MultLoop_and_154_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_601_rgt
      , and_dcpl_467});
  assign nand_198_cse = ~((fsm_output[3]) & (fsm_output[7]));
  assign and_472_m1c = or_dcpl_394 & IndexLoop_stage_0_2;
  assign and_471_rgt = and_dcpl_263 & and_dcpl_197 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_281_rgt
      = ((~ or_dcpl_584) & and_472_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_636_cse;
  assign MultLoop_and_152_rgt = or_dcpl_584 & and_472_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_108_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_788_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_474_m1c = or_dcpl_392 & IndexLoop_stage_0_2;
  assign or_1398_cse = (fsm_output[6:5]!=2'b00);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_250_rgt
      = (and_dcpl_255 & and_dcpl_261 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_607_cse;
  assign MultLoop_and_149_rgt = (~ or_dcpl_583) & and_474_m1c & and_dcpl_65;
  assign MultLoop_and_150_rgt = or_dcpl_583 & and_474_m1c & and_dcpl_65;
  assign and_476_m1c = or_dcpl_390 & IndexLoop_stage_0_2;
  assign and_475_rgt = and_dcpl_274 & and_dcpl_223 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_280_rgt
      = ((~ or_dcpl_582) & and_476_m1c & and_dcpl_65) | (and_dcpl_219 & and_dcpl_204
      & and_dcpl_60);
  assign MultLoop_and_148_rgt = or_dcpl_582 & and_476_m1c & and_dcpl_65;
  assign and_478_rgt = or_dcpl_518 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_110_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_802_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_480_m1c = or_dcpl_389 & IndexLoop_stage_0_2;
  assign or_1213_cse = (~ (fsm_output[5])) | (fsm_output[7]);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_249_rgt
      = (and_dcpl_266 & and_dcpl_235 & and_dcpl_65) | (and_dcpl_283 & and_dcpl_216
      & and_dcpl_60);
  assign MultLoop_and_145_rgt = (~ or_dcpl_581) & and_480_m1c & and_dcpl_65;
  assign MultLoop_and_146_rgt = or_dcpl_581 & and_480_m1c & and_dcpl_65;
  assign and_482_rgt = or_dcpl_520 & and_dcpl_176 & and_dcpl_60;
  assign nor_952_cse = ~((fsm_output[3]) | (fsm_output[4]) | (fsm_output[7]));
  assign or_1800_cse = (fsm_output[6]) | (fsm_output[2]);
  assign and_484_m1c = or_dcpl_388 & IndexLoop_stage_0_2;
  assign and_483_rgt = and_dcpl_263 & and_dcpl_223 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_279_rgt
      = ((~ or_dcpl_580) & and_484_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_539_cse;
  assign MultLoop_and_144_rgt = or_dcpl_580 & and_484_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_112_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_815_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_486_m1c = or_dcpl_386 & IndexLoop_stage_0_2;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_248_rgt
      = (and_dcpl_255 & and_dcpl_235 & and_dcpl_65) | (and_dcpl_486 & and_dcpl_204
      & and_dcpl_60);
  assign MultLoop_and_141_rgt = (~ or_dcpl_579) & and_486_m1c & and_dcpl_65;
  assign MultLoop_and_142_rgt = or_dcpl_579 & and_486_m1c & and_dcpl_65;
  assign and_489_rgt = or_dcpl_526 & and_dcpl_176 & and_dcpl_60;
  assign and_491_m1c = or_dcpl_384 & IndexLoop_stage_0_2;
  assign and_490_rgt = and_dcpl_247 & and_dcpl_197 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_278_rgt
      = ((~ or_dcpl_578) & and_491_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_439_cse;
  assign MultLoop_and_140_rgt = or_dcpl_578 & and_491_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_114_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_832_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_493_m1c = or_dcpl_383 & IndexLoop_stage_0_2;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_247_rgt
      = (and_dcpl_212 & and_dcpl_261 & and_dcpl_65) | (and_dcpl_486 & and_dcpl_216
      & and_dcpl_60);
  assign MultLoop_and_137_rgt = (~ or_dcpl_577) & and_493_m1c & and_dcpl_65;
  assign MultLoop_and_138_rgt = or_dcpl_577 & and_493_m1c & and_dcpl_65;
  assign and_495_rgt = or_dcpl_517 & and_dcpl_176 & and_dcpl_60;
  assign and_497_m1c = or_dcpl_382 & IndexLoop_stage_0_2;
  assign and_496_rgt = and_dcpl_181 & and_dcpl_197 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_396_cse
      = and_dcpl_415 & and_dcpl_216 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_277_rgt
      = ((~ or_dcpl_576) & and_497_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_396_cse;
  assign MultLoop_and_136_rgt = or_dcpl_576 & and_497_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_397_rgt
      = or_dcpl_558 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_116_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_846_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_501_m1c = or_dcpl_377 & IndexLoop_stage_0_2;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_246_rgt
      = (and_dcpl_200 & and_dcpl_261 & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_396_cse;
  assign MultLoop_and_133_rgt = (~ or_dcpl_575) & and_501_m1c & and_dcpl_65;
  assign MultLoop_and_134_rgt = or_dcpl_575 & and_501_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_117_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_850_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_503_m1c = or_dcpl_372 & IndexLoop_stage_0_2;
  assign and_502_rgt = and_dcpl_247 & and_dcpl_223 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_276_rgt
      = ((~ or_dcpl_574) & and_503_m1c & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_479_cse;
  assign MultLoop_and_132_rgt = or_dcpl_574 & and_503_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_118_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_856_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_505_m1c = or_dcpl_366 & IndexLoop_stage_0_2;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_245_rgt
      = (and_dcpl_212 & and_dcpl_235 & and_dcpl_65) | (and_dcpl_251 & and_dcpl_216
      & and_dcpl_60);
  assign MultLoop_and_129_rgt = (~ or_dcpl_573) & and_505_m1c & and_dcpl_65;
  assign MultLoop_and_130_rgt = or_dcpl_573 & and_505_m1c & and_dcpl_65;
  assign and_507_rgt = or_dcpl_559 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_119_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_862_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_509_m1c = or_dcpl_490 & IndexLoop_stage_0_2;
  assign and_508_rgt = and_dcpl_181 & and_dcpl_223 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_275_rgt
      = ((~ or_dcpl_572) & and_509_m1c & and_dcpl_65) | (and_dcpl_509 & and_dcpl_216
      & and_dcpl_60);
  assign MultLoop_and_128_rgt = or_dcpl_572 & and_509_m1c & and_dcpl_65;
  assign and_512_rgt = or_dcpl_495 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_120_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_867_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign and_514_m1c = or_dcpl_560 & IndexLoop_stage_0_2;
  assign mux_249_cse = MUX_s_1_2_2(or_864_cse, (fsm_output[7]), fsm_output[5]);
  assign and_513_rgt = and_dcpl_200 & and_dcpl_235 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_274_rgt
      = ((~ or_dcpl_571) & and_514_m1c & and_dcpl_65) | (and_dcpl_509 & and_dcpl_204
      & and_dcpl_60);
  assign MultLoop_and_126_rgt = or_dcpl_571 & and_514_m1c & and_dcpl_65;
  assign and_516_rgt = or_dcpl_561 & and_dcpl_176 & and_dcpl_60;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_121_ssc
      = core_wen & (and_dcpl_65 | and_dcpl_60 | (~ mux_872_itm)) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse;
  assign MultLoop_2_nor_m1c = ~((ROM_1i9_1o3_2fa806bf16b3e0d54016201674d036b62f_1!=3'b000));
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_371_m1c
      = or_dcpl_448 & (~ or_1479_cse);
  assign or_1298_cse = (~ (fsm_output[2])) | (fsm_output[6]) | (~ (fsm_output[7]));
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_129_cse
      = or_dcpl_559 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_63_nl
      = ~(or_dcpl_447 | or_1479_cse);
  assign MultLoop_and_253_nl = (~ or_dcpl_572) & or_dcpl_447 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_185_nl =
      or_dcpl_572 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_63_nl
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, ({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_1_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_2_reg}),
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_63_nl)
      , (MultLoop_and_253_nl) , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_185_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_62_nl
      = ~(or_dcpl_448 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_372_nl
      = (~ or_dcpl_571) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_371_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_184_nl =
      (or_dcpl_571 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_371_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_62_nl
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, ({reg_MultLoop_1_mux_64_itm_1_reg ,
      reg_MultLoop_1_mux_64_itm_1_1_reg}), {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_62_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_372_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_184_nl)});
  assign MultLoop_mux_129_nl = MUX_v_18_64_2((nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_63_nl),
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_1_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_6_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_8_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_9_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_10_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_58_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_59_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_60_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_61_1_sva_1_mx2,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_sva_1_mx2,
      (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_62_nl),
      IndexLoop_mux_1_tmp);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_30_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_32_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_128_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_29_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_33_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_96_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_28_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_34_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_97_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_27_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_35_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_98_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_26_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_36_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_99_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_25_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_37_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_100_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_24_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_38_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_101_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_23_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_39_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_102_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_22_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_40_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_103_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_21_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_41_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_104_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_20_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_42_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_105_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_19_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_43_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_106_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_18_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_44_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_107_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_17_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_45_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_108_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_16_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_46_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_109_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_15_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_47_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_110_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_14_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_48_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_111_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_13_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_49_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_112_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_12_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_50_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_113_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_11_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_51_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_114_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_10_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_52_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_115_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_9_nl =
      MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_53_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_116_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_8_nl =
      MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_54_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_117_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_7_nl =
      MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_55_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_118_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_6_nl =
      MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_56_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_119_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_5_nl =
      MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_57_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_120_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_4_nl =
      MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_58_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_121_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_3_nl =
      MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_59_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_122_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_2_nl =
      MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_60_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_123_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_1_nl =
      MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_61_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_124_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_nl = MUX_v_18_2_2(z_out_21,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_62_sva_1, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_125_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_63_nl
      = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_63_sva,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_129_cse);
  assign MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_nl
      = MUX_v_18_32_2((nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_30_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_29_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_28_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_27_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_26_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_25_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_24_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_23_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_22_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_21_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_20_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_19_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_18_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_17_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_16_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_15_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_14_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_13_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_12_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_11_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_10_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_9_nl), (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_8_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_7_nl), (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_6_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_5_nl), (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_4_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_3_nl), (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_2_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_1_nl), (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_63_nl),
      ROM_1i11_1o5_b94ddd86102738ded3ce1c444a799cda31_1);
  assign MultLoop_or_7_nl = (and_dcpl_65 & and_dcpl_424 & and_dcpl_325) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_465_cse;
  assign MultLoop_or_8_nl = ((~ or_dcpl_592) & MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_mx0c2)
      | ((((~ or_1420_tmp) & MultLoop_2_and_26_m1c) | (nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_11_cse
      & MultLoop_2_and_28_m1c) | (and_dcpl_176 & MultLoop_2_and_6_itm_1) | (nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_10_cse
      & MultLoop_2_and_29_m1c) | (nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_9_cse
      & MultLoop_2_and_30_m1c) | ((~ nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_or_8_cse)
      & MultLoop_2_and_31_m1c)) & and_dcpl_55);
  assign MultLoop_and_250_nl = or_dcpl_592 & MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_mx0c2;
  assign and_541_nl = or_dcpl_552 & and_dcpl_75 & and_dcpl_449;
  assign MultLoop_and_261_nl = ((or_1420_tmp & MultLoop_2_and_26_m1c) | (or_1479_cse
      & MultLoop_2_nor_m1c & IndexLoop_stage_0)) & and_dcpl_55;
  assign MultLoop_2_and_32_nl = (~ nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_11_cse)
      & MultLoop_2_and_28_m1c & and_dcpl_55;
  assign MultLoop_and_262_nl = (((~ nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_10_cse)
      & MultLoop_2_and_29_m1c) | (and_dcpl_176 & (~ MultLoop_2_and_6_itm_1))) & and_dcpl_55;
  assign MultLoop_2_and_37_nl = (~ nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_9_cse)
      & MultLoop_2_and_30_m1c & and_dcpl_55;
  assign MultLoop_2_and_39_nl = nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_or_8_cse
      & MultLoop_2_and_31_m1c & and_dcpl_55;
  assign mux_891_nl = MUX_s_1_2_2(nor_942_cse, mux_456_cse, fsm_output[1]);
  assign mux_892_nl = MUX_s_1_2_2(nor_310_cse, (mux_891_nl), fsm_output[0]);
  assign and_542_nl = (~ (mux_892_nl)) & and_dcpl_100;
  assign MultLoop_mux1h_60_rgt = MUX1HOT_v_18_12_2((MultLoop_mux_129_nl), z_out_20,
      z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_10_1_sva_1,
      (MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_nl),
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_11_sva_1, ({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_1_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_2_reg}),
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_1_sva_1, nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_2_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_3_sva_1, nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_4_sva_1,
      ({6'b000000 , CALC_SOFTMAX_LOOP_6_or_cse}), {and_dcpl_82 , (MultLoop_or_7_nl)
      , (MultLoop_or_8_nl) , (MultLoop_and_250_nl) , and_dcpl_77 , (and_541_nl) ,
      (MultLoop_and_261_nl) , (MultLoop_2_and_32_nl) , (MultLoop_and_262_nl) , (MultLoop_2_and_37_nl)
      , (MultLoop_2_and_39_nl) , (and_542_nl)});
  assign and_2630_cse = ((ROM_1i9_1o3_2fa806bf16b3e0d54016201674d036b62f_1[1:0]!=2'b00))
      & (ROM_1i9_1o3_2fa806bf16b3e0d54016201674d036b62f_1[2]);
  assign and_2631_cse = (fsm_output[7]) & (fsm_output[4]);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_128_cse
      = or_dcpl_561 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_62_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_0_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_128_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_31_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_1_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_96_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_32_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_2_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_97_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_33_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_3_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_98_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_34_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_4_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_99_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_35_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_5_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_100_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_36_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_6_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_101_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_37_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_7_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_102_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_38_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_8_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_103_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_39_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_9_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_104_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_40_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_10_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_105_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_41_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_11_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_106_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_42_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_12_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_107_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_43_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_13_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_108_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_44_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_14_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_109_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_45_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_15_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_110_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_46_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_16_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_111_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_47_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_17_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_112_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_48_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_18_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_113_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_49_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_19_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_114_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_50_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_20_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_115_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_51_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_21_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_116_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_52_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_22_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_117_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_53_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_23_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_118_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_54_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_24_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_119_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_55_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_25_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_120_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_56_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_26_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_121_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_57_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_27_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_122_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_58_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_28_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_123_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_59_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_29_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_124_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_60_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_30_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_125_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_61_nl
      = MUX_v_18_2_2(z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_31_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_129_cse);
  assign MultLoop_1_mux_64_nl = MUX_v_18_32_2((nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_62_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_31_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_32_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_33_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_34_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_35_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_36_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_37_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_38_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_39_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_40_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_41_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_42_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_43_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_44_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_45_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_46_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_47_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_48_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_49_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_50_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_51_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_52_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_53_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_54_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_55_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_56_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_57_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_58_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_59_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_60_nl),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_mux_61_nl),
      ROM_1i11_1o5_b94ddd86102738ded3ce1c444a799cda31_1);
  assign MultLoop_1_or_3_nl = (((and_dcpl_247 & and_dcpl_178) | ((~ or_dcpl_448)
      & and_dcpl_185)) & and_dcpl_65) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_456_cse
      | (((nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_15_cse
      & MultLoop_2_and_20_m1c) | ((~ or_1419_tmp) & MultLoop_2_and_21_m1c) | (nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_14_cse
      & MultLoop_2_and_25_m1c) | (nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_13_cse
      & MultLoop_2_and_24_m1c) | ((~ nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_or_9_cse)
      & MultLoop_2_and_23_m1c)) & and_dcpl_55);
  assign MultLoop_1_or_4_nl = ((((~ or_dcpl_574) & and_550_m1c) | ((~ or_dcpl_571)
      & or_dcpl_448 & and_dcpl_185)) & and_dcpl_65) | (and_dcpl_176 & MultLoop_2_and_7_itm_1
      & and_dcpl_55);
  assign MultLoop_and_247_nl = or_dcpl_574 & and_550_m1c & and_dcpl_65;
  assign and_547_nl = or_dcpl_554 & and_dcpl_75 & and_dcpl_449;
  assign MultLoop_2_and_42_nl = (~ nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_15_cse)
      & MultLoop_2_and_20_m1c & and_dcpl_55;
  assign MultLoop_1_and_66_nl = ((or_1419_tmp & MultLoop_2_and_21_m1c) | (or_1479_cse
      & MultLoop_2_and_m1c & IndexLoop_stage_0)) & and_dcpl_55;
  assign MultLoop_2_and_51_nl = nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_or_9_cse
      & MultLoop_2_and_23_m1c & and_dcpl_55;
  assign MultLoop_2_and_47_nl = (~ nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_13_cse)
      & MultLoop_2_and_24_m1c & and_dcpl_55;
  assign MultLoop_2_and_45_nl = (~ nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_14_cse)
      & MultLoop_2_and_25_m1c & and_dcpl_55;
  assign and_552_nl = and_dcpl_176 & (~ MultLoop_2_and_7_itm_1) & and_dcpl_55;
  assign mux_460_nl = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), and_817_cse);
  assign mux_901_nl = MUX_s_1_2_2(nor_310_cse, (mux_460_nl), fsm_output[0]);
  assign and_548_nl = (~ (mux_901_nl)) & and_dcpl_100;
  assign MultLoop_1_mux1h_65_rgt = MUX1HOT_v_18_13_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
      z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_1_1_sva_1,
      (MultLoop_1_mux_64_nl), nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_10_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_8_sva_1, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2,
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_5_sva_1, nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_6_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_7_sva_1, nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_1_sva_1,
      ({6'b000000 , CALC_SOFTMAX_LOOP_6_or_cse}), {and_dcpl_155 , (MultLoop_1_or_3_nl)
      , (MultLoop_1_or_4_nl) , (MultLoop_and_247_nl) , and_dcpl_77 , (and_547_nl)
      , (MultLoop_2_and_42_nl) , (MultLoop_1_and_66_nl) , (MultLoop_2_and_51_nl)
      , (MultLoop_2_and_47_nl) , (MultLoop_2_and_45_nl) , (and_552_nl) , (and_548_nl)});
  assign nand_191_cse = ~((InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b11111) & (~
      IndexLoop_asn_3_itm_1));
  assign nor_560_cse = ~((MultLoop_2_1_acc_3_tmp[1:0]!=2'b00));
  assign and_554_m1c = or_dcpl_431 & IndexLoop_stage_0_2;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_62_cse
      = core_wen & (and_dcpl_65 | and_dcpl_158 | and_dcpl_60);
  assign or_1393_nl = IndexLoop_stage_0 | (~ or_dcpl_561);
  assign nor_215_nl = ~(IndexLoop_stage_0 | (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1!=5'b00000));
  assign mux_907_nl = MUX_s_1_2_2((or_1393_nl), (nor_215_nl), IndexLoop_asn_3_itm_1);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_126_tmp
      = (or_dcpl_561 & and_dcpl_185) | (~((mux_907_nl) & IndexLoop_stage_0_2));
  assign and_556_m1c = or_dcpl_429 & IndexLoop_stage_0_2;
  assign or_1392_nl = IndexLoop_stage_0 | ((nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1==5'b11111));
  assign nor_214_nl = ~(IndexLoop_stage_0 | or_dcpl_559);
  assign mux_908_nl = MUX_s_1_2_2((or_1392_nl), (nor_214_nl), IndexLoop_asn_3_itm_1);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_127_tmp
      = (or_dcpl_559 & and_dcpl_185) | (~((mux_908_nl) & IndexLoop_stage_0_2));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_cse_16_15
      = MUX_v_2_2_2(2'b00, (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg[1:0]),
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_cse_14_12
      = MUX_v_3_2_2(3'b000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_1_reg,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_cse_11_0
      = MUX_v_12_2_2(12'b000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_2_reg,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer4_t_layer5_t_relu_config5_for_nnet_relu_layer4_t_layer5_t_relu_config5_for_and_cse
      = MUX_v_17_2_2(17'b00000000000000000, (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_0_sva_1[16:0]),
      (z_out_23_22_8[10]));
  assign and_558_ssc = and_dcpl_59 & and_dcpl_159;
  assign nor_554_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[4]));
  assign nor_555_nl = ~((fsm_output[7]) | (fsm_output[6]) | (fsm_output[4]));
  assign nor_556_nl = ~((~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[4])));
  assign mux_1242_nl = MUX_s_1_2_2((nor_555_nl), (nor_556_nl), fsm_output[2]);
  assign mux_1243_cse = MUX_s_1_2_2((nor_554_nl), (mux_1242_nl), fsm_output[0]);
  assign and_2623_nl = (fsm_output[1]) & mux_1243_cse;
  assign nor_557_nl = ~(and_2642_cse | (~ (fsm_output[7])) | (fsm_output[6]) | (~
      (fsm_output[4])));
  assign mux_1244_nl = MUX_s_1_2_2((and_2623_nl), (nor_557_nl), fsm_output[3]);
  assign and_2617_ssc = (mux_1244_nl) & (~ (fsm_output[5])) & core_wen;
  assign and_566_rgt = and_dcpl_59 & and_dcpl_51;
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_2_ssc = core_wen & mux_tmp_911;
  assign and_568_rgt = and_dcpl_59 & and_dcpl_519;
  assign mux_927_nl = MUX_s_1_2_2(mux_tmp_926, mux_tmp_911, fsm_output[0]);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_3_ssc = core_wen & (mux_927_nl);
  assign MultLoop_2_and_5_itm = (ROM_1i9_1o3_2fa806bf16b3e0d54016201674d036b62f_1==3'b011);
  assign MultLoop_2_and_6_itm = (ROM_1i9_1o3_2fa806bf16b3e0d54016201674d036b62f_1==3'b010);
  assign MultLoop_2_and_7_itm = (ROM_1i9_1o3_2fa806bf16b3e0d54016201674d036b62f_1==3'b001);
  assign MultLoop_2_and_cse = core_wen & (and_dcpl_55 | and_dcpl_520);
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_10_18_6_true_AC_TRN_AC_SAT_18_2_AC_TRN_AC_SAT_exp_arr_and_cse
      = core_wen & (~(or_dcpl_455 | or_dcpl_607 | or_1875_cse));
  assign operator_67_47_false_AC_TRN_AC_WRAP_and_1_cse = core_wen & (~(or_dcpl_455
      | or_dcpl_607 | or_dcpl_465));
  assign and_727_nl = and_dcpl_100 & and_dcpl_154;
  assign SUM_EXP_LOOP_mux_1_rgt = MUX_v_70_2_2(({2'b00 , (z_out_24[67:0])}), (z_out_10[69:0]),
      and_727_nl);
  assign operator_67_47_false_AC_TRN_AC_WRAP_and_5_cse = core_wen & (~(or_dcpl_455
      | or_dcpl_467));
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_245_m1c
      = or_dcpl_446 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_nl
      = ~(or_dcpl_446 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_368_nl
      = (~ or_dcpl_573) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_245_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_183_nl =
      (or_dcpl_573 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_245_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_368_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_183_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_243_m1c
      = or_dcpl_445 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_1_nl
      = ~(or_dcpl_445 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_366_nl
      = (~ or_dcpl_574) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_243_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_182_nl =
      (or_dcpl_574 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_243_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_1_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_1_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_1_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_366_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_182_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_241_m1c
      = or_dcpl_444 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_2_nl
      = ~(or_dcpl_444 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_364_nl
      = (~ or_dcpl_575) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_241_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_181_nl =
      (or_dcpl_575 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_241_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_61_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_61_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_2_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_364_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_181_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_239_m1c
      = or_dcpl_443 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_3_nl
      = ~(or_dcpl_443 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_362_nl
      = (~ or_dcpl_576) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_239_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_180_nl =
      (or_dcpl_576 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_239_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_3_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_362_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_180_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_237_m1c
      = or_dcpl_442 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_4_nl
      = ~(or_dcpl_442 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_360_nl
      = (~ or_dcpl_577) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_237_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_179_nl =
      (or_dcpl_577 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_237_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_60_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_60_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_4_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_360_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_179_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_235_m1c
      = or_dcpl_441 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_5_nl
      = ~(or_dcpl_441 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_358_nl
      = (~ or_dcpl_578) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_235_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_178_nl =
      (or_dcpl_578 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_235_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_5_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_358_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_178_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_233_m1c
      = or_dcpl_440 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_6_nl
      = ~(or_dcpl_440 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_356_nl
      = (~ or_dcpl_579) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_233_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_177_nl =
      (or_dcpl_579 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_233_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_59_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_59_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_6_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_356_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_177_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_231_m1c
      = or_dcpl_439 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_7_nl
      = ~(or_dcpl_439 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_354_nl
      = (~ or_dcpl_580) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_231_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_176_nl =
      (or_dcpl_580 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_231_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_7_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_354_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_176_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_229_m1c
      = or_dcpl_438 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_8_nl
      = ~(or_dcpl_438 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_352_nl
      = (~ or_dcpl_581) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_229_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_175_nl =
      (or_dcpl_581 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_229_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_58_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_58_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_8_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_352_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_175_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_227_m1c
      = or_dcpl_437 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_9_nl
      = ~(or_dcpl_437 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_350_nl
      = (~ or_dcpl_582) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_227_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_174_nl =
      (or_dcpl_582 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_227_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_9_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_350_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_174_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_225_m1c
      = or_dcpl_436 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_10_nl
      = ~(or_dcpl_436 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_348_nl
      = (~ or_dcpl_583) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_225_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_173_nl =
      (or_dcpl_583 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_225_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_10_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_348_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_173_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_223_m1c
      = or_dcpl_435 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_11_nl
      = ~(or_dcpl_435 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_346_nl
      = (~ or_dcpl_584) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_223_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_172_nl =
      (or_dcpl_584 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_223_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_6_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_6_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_11_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_346_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_172_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_221_m1c
      = or_dcpl_434 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_12_nl
      = ~(or_dcpl_434 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_344_nl
      = (~ or_dcpl_585) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_221_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_171_nl =
      (or_dcpl_585 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_221_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_12_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_344_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_171_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_219_m1c
      = or_dcpl_433 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_13_nl
      = ~(or_dcpl_433 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_342_nl
      = (~ or_dcpl_586) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_219_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_170_nl =
      (or_dcpl_586 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_219_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_13_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_342_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_170_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_217_m1c
      = or_dcpl_432 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_14_nl
      = ~(or_dcpl_432 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_340_nl
      = (~ or_dcpl_587) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_217_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_169_nl =
      (or_dcpl_587 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_217_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_14_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_340_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_169_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_215_m1c
      = or_dcpl_431 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_15_nl
      = ~(or_dcpl_431 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_338_nl
      = (~ or_dcpl_588) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_215_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_168_nl =
      (or_dcpl_588 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_215_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_8_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_8_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_15_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_338_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_168_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_213_m1c
      = or_dcpl_430 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_16_nl
      = ~(or_dcpl_430 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_336_nl
      = (~ or_dcpl_589) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_213_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_167_nl =
      (or_dcpl_589 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_213_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_16_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_336_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_167_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_211_m1c
      = or_dcpl_429 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_17_nl
      = ~(or_dcpl_429 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_334_nl
      = (~ or_dcpl_590) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_211_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_166_nl =
      (or_dcpl_590 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_211_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_9_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_9_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_17_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_334_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_166_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_209_m1c
      = or_dcpl_428 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_18_nl
      = ~(or_dcpl_428 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_332_nl
      = (~ or_dcpl_591) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_209_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_165_nl =
      (or_dcpl_591 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_209_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_18_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_332_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_165_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_207_m1c
      = or_dcpl_427 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_19_nl
      = ~(or_dcpl_427 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_330_nl
      = (~ or_dcpl_592) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_207_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_164_nl =
      (or_dcpl_592 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_207_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_10_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_10_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_19_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_330_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_164_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_205_m1c
      = or_dcpl_426 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_20_nl
      = ~(or_dcpl_426 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_328_nl
      = (~ or_dcpl_593) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_205_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_163_nl =
      (or_dcpl_593 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_205_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_20_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_328_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_163_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_203_m1c
      = or_dcpl_425 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_21_nl
      = ~(or_dcpl_425 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_326_nl
      = (~ or_dcpl_594) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_203_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_162_nl =
      (or_dcpl_594 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_203_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_21_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_326_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_162_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_201_m1c
      = or_dcpl_424 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_22_nl
      = ~(or_dcpl_424 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_324_nl
      = (~ or_dcpl_595) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_201_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_161_nl =
      (or_dcpl_595 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_201_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_22_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_324_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_161_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_199_m1c
      = or_dcpl_423 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_23_nl
      = ~(or_dcpl_423 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_322_nl
      = (~ or_dcpl_596) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_199_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_160_nl =
      (or_dcpl_596 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_199_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_23_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_322_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_160_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_197_m1c
      = or_dcpl_422 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_24_nl
      = ~(or_dcpl_422 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_320_nl
      = (~ or_dcpl_597) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_197_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_159_nl =
      (or_dcpl_597 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_197_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_24_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_320_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_159_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_195_m1c
      = or_dcpl_421 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_25_nl
      = ~(or_dcpl_421 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_318_nl
      = (~ or_dcpl_598) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_195_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_158_nl =
      (or_dcpl_598 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_195_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_25_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_318_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_158_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_193_m1c
      = or_dcpl_420 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_26_nl
      = ~(or_dcpl_420 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_316_nl
      = (~ or_dcpl_599) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_193_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_157_nl =
      (or_dcpl_599 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_193_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_26_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_316_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_157_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_191_m1c
      = or_dcpl_419 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_27_nl
      = ~(or_dcpl_419 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_314_nl
      = (~ or_dcpl_600) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_191_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_156_nl =
      (or_dcpl_600 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_191_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_27_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_314_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_156_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_189_m1c
      = or_dcpl_418 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_28_nl
      = ~(or_dcpl_418 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_312_nl
      = (~ or_dcpl_601) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_189_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_155_nl =
      (or_dcpl_601 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_189_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_28_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_312_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_155_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_187_m1c
      = or_dcpl_417 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_29_nl
      = ~(or_dcpl_417 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_310_nl
      = (~ or_dcpl_602) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_187_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_154_nl =
      (or_dcpl_602 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_187_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_29_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_310_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_154_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_185_m1c
      = or_dcpl_416 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_30_nl
      = ~(or_dcpl_416 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_308_nl
      = (~ or_dcpl_602) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_185_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_153_nl =
      (or_dcpl_602 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_185_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_30_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_308_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_153_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_183_m1c
      = or_dcpl_415 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_31_nl
      = ~(or_dcpl_415 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_306_nl
      = (~ or_dcpl_601) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_183_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_152_nl =
      (or_dcpl_601 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_183_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_31_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_306_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_152_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_181_m1c
      = or_dcpl_414 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_32_nl
      = ~(or_dcpl_414 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_304_nl
      = (~ or_dcpl_600) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_181_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_151_nl =
      (or_dcpl_600 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_181_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_32_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_304_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_151_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_179_m1c
      = or_dcpl_413 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_33_nl
      = ~(or_dcpl_413 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_302_nl
      = (~ or_dcpl_599) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_179_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_150_nl =
      (or_dcpl_599 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_179_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_33_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_302_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_150_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_177_m1c
      = or_dcpl_412 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_34_nl
      = ~(or_dcpl_412 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_300_nl
      = (~ or_dcpl_598) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_177_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_149_nl =
      (or_dcpl_598 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_177_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_34_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_300_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_149_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_175_m1c
      = or_dcpl_411 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_35_nl
      = ~(or_dcpl_411 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_298_nl
      = (~ or_dcpl_597) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_175_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_148_nl =
      (or_dcpl_597 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_175_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_35_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_298_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_148_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_173_m1c
      = or_dcpl_410 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_36_nl
      = ~(or_dcpl_410 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_296_nl
      = (~ or_dcpl_596) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_173_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_147_nl =
      (or_dcpl_596 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_173_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_36_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_296_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_147_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_171_m1c
      = or_dcpl_409 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_37_nl
      = ~(or_dcpl_409 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_294_nl
      = (~ or_dcpl_595) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_171_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_146_nl =
      (or_dcpl_595 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_171_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_37_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_294_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_146_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_169_m1c
      = or_dcpl_408 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_38_nl
      = ~(or_dcpl_408 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_292_nl
      = (~ or_dcpl_594) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_169_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_145_nl =
      (or_dcpl_594 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_169_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_38_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_292_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_145_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_167_m1c
      = or_dcpl_407 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_39_nl
      = ~(or_dcpl_407 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_290_nl
      = (~ or_dcpl_593) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_167_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_144_nl =
      (or_dcpl_593 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_167_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_39_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_290_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_144_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_165_m1c
      = or_dcpl_406 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_40_nl
      = ~(or_dcpl_406 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_288_nl
      = (~ or_dcpl_592) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_165_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_143_nl =
      (or_dcpl_592 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_165_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_40_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_288_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_143_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_163_m1c
      = or_dcpl_405 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_41_nl
      = ~(or_dcpl_405 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_286_nl
      = (~ or_dcpl_591) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_163_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_142_nl =
      (or_dcpl_591 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_163_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_41_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_286_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_142_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_161_m1c
      = or_dcpl_404 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_42_nl
      = ~(or_dcpl_404 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_284_nl
      = (~ or_dcpl_590) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_161_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_141_nl =
      (or_dcpl_590 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_161_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_42_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_284_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_141_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_159_m1c
      = or_dcpl_402 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_43_nl
      = ~(or_dcpl_402 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_282_nl
      = (~ or_dcpl_589) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_159_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_140_nl =
      (or_dcpl_589 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_159_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_43_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_282_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_140_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_157_m1c
      = or_dcpl_400 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_44_nl
      = ~(or_dcpl_400 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_280_nl
      = (~ or_dcpl_588) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_157_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_139_nl =
      (or_dcpl_588 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_157_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_44_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_280_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_139_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_155_m1c
      = or_dcpl_398 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_45_nl
      = ~(or_dcpl_398 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_278_nl
      = (~ or_dcpl_587) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_155_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_138_nl =
      (or_dcpl_587 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_155_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_45_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_278_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_138_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_153_m1c
      = or_dcpl_396 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_46_nl
      = ~(or_dcpl_396 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_276_nl
      = (~ or_dcpl_586) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_153_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_137_nl =
      (or_dcpl_586 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_153_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_46_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_276_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_137_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_151_m1c
      = or_dcpl_395 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_47_nl
      = ~(or_dcpl_395 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_274_nl
      = (~ or_dcpl_585) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_151_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_136_nl =
      (or_dcpl_585 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_151_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_47_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_274_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_136_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_149_m1c
      = or_dcpl_394 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_48_nl
      = ~(or_dcpl_394 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_272_nl
      = (~ or_dcpl_584) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_149_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_135_nl =
      (or_dcpl_584 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_149_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_48_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_272_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_135_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_147_m1c
      = or_dcpl_392 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_49_nl
      = ~(or_dcpl_392 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_270_nl
      = (~ or_dcpl_583) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_147_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_134_nl =
      (or_dcpl_583 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_147_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_49_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_270_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_134_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_145_m1c
      = or_dcpl_390 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_50_nl
      = ~(or_dcpl_390 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_268_nl
      = (~ or_dcpl_582) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_145_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_133_nl =
      (or_dcpl_582 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_145_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_50_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_268_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_133_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_143_m1c
      = or_dcpl_389 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_51_nl
      = ~(or_dcpl_389 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_266_nl
      = (~ or_dcpl_581) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_143_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_132_nl =
      (or_dcpl_581 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_143_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_51_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_266_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_132_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_141_m1c
      = or_dcpl_388 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_52_nl
      = ~(or_dcpl_388 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_264_nl
      = (~ or_dcpl_580) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_141_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_131_nl =
      (or_dcpl_580 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_141_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_52_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_264_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_131_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_139_m1c
      = or_dcpl_386 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_53_nl
      = ~(or_dcpl_386 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_262_nl
      = (~ or_dcpl_579) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_139_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_130_nl =
      (or_dcpl_579 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_139_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_53_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_262_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_130_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_137_m1c
      = or_dcpl_384 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_54_nl
      = ~(or_dcpl_384 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_260_nl
      = (~ or_dcpl_578) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_137_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_129_nl =
      (or_dcpl_578 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_137_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_54_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_260_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_129_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_135_m1c
      = or_dcpl_383 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_55_nl
      = ~(or_dcpl_383 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_258_nl
      = (~ or_dcpl_577) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_135_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_128_nl =
      (or_dcpl_577 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_135_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_55_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_258_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_128_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_133_m1c
      = or_dcpl_382 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_56_nl
      = ~(or_dcpl_382 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_256_nl
      = (~ or_dcpl_576) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_133_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_127_nl =
      (or_dcpl_576 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_133_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_56_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_256_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_127_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_131_m1c
      = or_dcpl_377 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_57_nl
      = ~(or_dcpl_377 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_254_nl
      = (~ or_dcpl_575) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_131_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_126_nl =
      (or_dcpl_575 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_131_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_57_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_254_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_126_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_129_m1c
      = or_dcpl_372 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_58_nl
      = ~(or_dcpl_372 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_252_nl
      = (~ or_dcpl_574) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_129_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_125_nl =
      (or_dcpl_574 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_129_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_58_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_252_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_125_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_127_m1c
      = or_dcpl_366 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_59_nl
      = ~(or_dcpl_366 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_250_nl
      = (~ or_dcpl_573) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_127_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_124_nl =
      (or_dcpl_573 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_127_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_59_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_250_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_124_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_125_m1c
      = or_dcpl_490 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_60_nl
      = ~(or_dcpl_490 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_248_nl
      = (~ or_dcpl_572) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_125_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_123_nl =
      (or_dcpl_572 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_125_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_60_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_248_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_123_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_123_m1c
      = or_dcpl_560 & (~ or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_61_nl
      = ~(or_dcpl_560 | or_1479_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_246_nl
      = (~ or_dcpl_571) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_123_m1c;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_122_nl =
      (or_dcpl_571 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_123_m1c)
      | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_sva_1_mx2
      = MUX1HOT_v_18_3_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_sva_1,
      {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_61_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_246_nl)
      , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_122_nl)});
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_125_cse
      = or_dcpl_513 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_124_cse
      = or_dcpl_517 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_123_cse
      = or_dcpl_526 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_122_cse
      = or_dcpl_520 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_121_cse
      = or_dcpl_525 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_120_cse
      = or_dcpl_528 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_119_cse
      = or_dcpl_531 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_118_cse
      = or_dcpl_533 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_117_cse
      = or_dcpl_534 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_116_cse
      = or_dcpl_535 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_115_cse
      = or_dcpl_516 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_114_cse
      = or_dcpl_541 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_113_cse
      = or_dcpl_522 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_112_cse
      = or_dcpl_547 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_111_cse
      = or_dcpl_548 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_110_cse
      = or_dcpl_546 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_109_cse
      = or_dcpl_543 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_108_cse
      = or_dcpl_538 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_107_cse
      = or_dcpl_537 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_106_cse
      = or_dcpl_552 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_105_cse
      = or_dcpl_554 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_104_cse
      = or_dcpl_529 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_103_cse
      = or_dcpl_501 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_102_cse
      = or_dcpl_505 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_101_cse
      = or_dcpl_518 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_100_cse
      = or_dcpl_545 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_99_cse
      = or_dcpl_556 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_98_cse
      = or_dcpl_558 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_97_cse
      = or_dcpl_551 | or_1479_cse;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_96_cse
      = or_dcpl_495 | or_1479_cse;
  assign IndexLoop_mux_1_tmp = MUX_v_6_16_2(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc15_sva,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc0_sva,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc1_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc2_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc3_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc4_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc5_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc6_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc7_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc8_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc9_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc10_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc11_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc12_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc13_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc14_sva_1,
      InitAccumLoop_2_iacc_3_0_sva);
  assign InitAccumLoop_2_slc_InitAccumLoop_2_asn_18_17_0_ctmp_sva_1 = MUX_v_18_10_2((b6_rsci_idat[17:0]),
      (b6_rsci_idat[35:18]), (b6_rsci_idat[53:36]), (b6_rsci_idat[71:54]), (b6_rsci_idat[89:72]),
      (b6_rsci_idat[107:90]), (b6_rsci_idat[125:108]), (b6_rsci_idat[143:126]), (b6_rsci_idat[161:144]),
      (b6_rsci_idat[179:162]), InitAccumLoop_2_iacc_3_0_sva);
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_2_nor_2_nl = ~(MUX_v_15_2_2(({(reg_MultLoop_1_mux_64_itm_1_reg[2:0])
      , reg_MultLoop_1_mux_64_itm_1_1_reg}), 15'b111111111111111, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_2_sva_mx0w1));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_2_and_nl = (reg_MultLoop_1_mux_64_itm_1_reg[5])
      & (~((reg_MultLoop_1_mux_64_itm_1_reg[4:3]==2'b11)));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_2_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl
      = ~(MUX_v_15_2_2((nnet_softmax_layer6_t_result_t_softmax_config7_for_2_nor_2_nl),
      15'b111111111111111, (nnet_softmax_layer6_t_result_t_softmax_config7_for_2_and_nl)));
  assign IndexLoop_ir_mux_nl = MUX_v_15_2_2((z_out_12[14:0]), (nnet_softmax_layer6_t_result_t_softmax_config7_for_2_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_nl),
      and_dcpl_520);
  assign or_12_nl = (fsm_output[1]) | nand_198_cse;
  assign or_1283_nl = (~ (fsm_output[1])) | (fsm_output[3]) | (fsm_output[7]);
  assign mux_884_nl = MUX_s_1_2_2((or_12_nl), (or_1283_nl), fsm_output[0]);
  assign nor_373_nl = ~((mux_884_nl) | or_1398_cse | (fsm_output[4]) | (fsm_output[2]));
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_3_14_0
      = MUX_v_15_2_2(15'b000000000000000, (IndexLoop_ir_mux_nl), (nor_373_nl));
  assign nl_IndexLoop_acc_nl = conv_u2s_6_7(z_out_13[14:9]) + 7'b1001111;
  assign IndexLoop_acc_nl = nl_IndexLoop_acc_nl[6:0];
  assign nl_ReuseLoop_acc_nl = conv_u2s_6_7(z_out_12[14:9]) + 7'b1001111;
  assign ReuseLoop_acc_nl = nl_ReuseLoop_acc_nl[6:0];
  assign IndexLoop_IndexLoop_nor_tmp = ~((readslicef_7_1_6((IndexLoop_acc_nl))) |
      (readslicef_7_1_6((ReuseLoop_acc_nl))));
  assign InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1
      = MUX_v_18_64_2((b2_rsci_idat[17:0]), (b2_rsci_idat[35:18]), (b2_rsci_idat[53:36]),
      (b2_rsci_idat[71:54]), (b2_rsci_idat[89:72]), (b2_rsci_idat[107:90]), (b2_rsci_idat[125:108]),
      (b2_rsci_idat[143:126]), (b2_rsci_idat[161:144]), (b2_rsci_idat[179:162]),
      (b2_rsci_idat[197:180]), (b2_rsci_idat[215:198]), (b2_rsci_idat[233:216]),
      (b2_rsci_idat[251:234]), (b2_rsci_idat[269:252]), (b2_rsci_idat[287:270]),
      (b2_rsci_idat[305:288]), (b2_rsci_idat[323:306]), (b2_rsci_idat[341:324]),
      (b2_rsci_idat[359:342]), (b2_rsci_idat[377:360]), (b2_rsci_idat[395:378]),
      (b2_rsci_idat[413:396]), (b2_rsci_idat[431:414]), (b2_rsci_idat[449:432]),
      (b2_rsci_idat[467:450]), (b2_rsci_idat[485:468]), (b2_rsci_idat[503:486]),
      (b2_rsci_idat[521:504]), (b2_rsci_idat[539:522]), (b2_rsci_idat[557:540]),
      (b2_rsci_idat[575:558]), (b2_rsci_idat[593:576]), (b2_rsci_idat[611:594]),
      (b2_rsci_idat[629:612]), (b2_rsci_idat[647:630]), (b2_rsci_idat[665:648]),
      (b2_rsci_idat[683:666]), (b2_rsci_idat[701:684]), (b2_rsci_idat[719:702]),
      (b2_rsci_idat[737:720]), (b2_rsci_idat[755:738]), (b2_rsci_idat[773:756]),
      (b2_rsci_idat[791:774]), (b2_rsci_idat[809:792]), (b2_rsci_idat[827:810]),
      (b2_rsci_idat[845:828]), (b2_rsci_idat[863:846]), (b2_rsci_idat[881:864]),
      (b2_rsci_idat[899:882]), (b2_rsci_idat[917:900]), (b2_rsci_idat[935:918]),
      (b2_rsci_idat[953:936]), (b2_rsci_idat[971:954]), (b2_rsci_idat[989:972]),
      (b2_rsci_idat[1007:990]), (b2_rsci_idat[1025:1008]), (b2_rsci_idat[1043:1026]),
      (b2_rsci_idat[1061:1044]), (b2_rsci_idat[1079:1062]), (b2_rsci_idat[1097:1080]),
      (b2_rsci_idat[1115:1098]), (b2_rsci_idat[1133:1116]), (b2_rsci_idat[1151:1134]),
      InitAccumLoop_1_iacc_6_0_sva_5_0);
  assign InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1
      = MUX_v_18_64_2((b4_rsci_idat[17:0]), (b4_rsci_idat[35:18]), (b4_rsci_idat[53:36]),
      (b4_rsci_idat[71:54]), (b4_rsci_idat[89:72]), (b4_rsci_idat[107:90]), (b4_rsci_idat[125:108]),
      (b4_rsci_idat[143:126]), (b4_rsci_idat[161:144]), (b4_rsci_idat[179:162]),
      (b4_rsci_idat[197:180]), (b4_rsci_idat[215:198]), (b4_rsci_idat[233:216]),
      (b4_rsci_idat[251:234]), (b4_rsci_idat[269:252]), (b4_rsci_idat[287:270]),
      (b4_rsci_idat[305:288]), (b4_rsci_idat[323:306]), (b4_rsci_idat[341:324]),
      (b4_rsci_idat[359:342]), (b4_rsci_idat[377:360]), (b4_rsci_idat[395:378]),
      (b4_rsci_idat[413:396]), (b4_rsci_idat[431:414]), (b4_rsci_idat[449:432]),
      (b4_rsci_idat[467:450]), (b4_rsci_idat[485:468]), (b4_rsci_idat[503:486]),
      (b4_rsci_idat[521:504]), (b4_rsci_idat[539:522]), (b4_rsci_idat[557:540]),
      (b4_rsci_idat[575:558]), (b4_rsci_idat[593:576]), (b4_rsci_idat[611:594]),
      (b4_rsci_idat[629:612]), (b4_rsci_idat[647:630]), (b4_rsci_idat[665:648]),
      (b4_rsci_idat[683:666]), (b4_rsci_idat[701:684]), (b4_rsci_idat[719:702]),
      (b4_rsci_idat[737:720]), (b4_rsci_idat[755:738]), (b4_rsci_idat[773:756]),
      (b4_rsci_idat[791:774]), (b4_rsci_idat[809:792]), (b4_rsci_idat[827:810]),
      (b4_rsci_idat[845:828]), (b4_rsci_idat[863:846]), (b4_rsci_idat[881:864]),
      (b4_rsci_idat[899:882]), (b4_rsci_idat[917:900]), (b4_rsci_idat[935:918]),
      (b4_rsci_idat[953:936]), (b4_rsci_idat[971:954]), (b4_rsci_idat[989:972]),
      (b4_rsci_idat[1007:990]), (b4_rsci_idat[1025:1008]), (b4_rsci_idat[1043:1026]),
      (b4_rsci_idat[1061:1044]), (b4_rsci_idat[1079:1062]), (b4_rsci_idat[1097:1080]),
      (b4_rsci_idat[1115:1098]), (b4_rsci_idat[1133:1116]), (b4_rsci_idat[1151:1134]),
      InitAccumLoop_1_iacc_6_0_sva_5_0);
  assign MultLoop_1_slc_input1_18_17_0_cse_sva_1 = MUX_v_18_784_2((input1_rsci_idat_mxwt[17:0]),
      (input1_rsci_idat_mxwt[35:18]), (input1_rsci_idat_mxwt[53:36]), (input1_rsci_idat_mxwt[71:54]),
      (input1_rsci_idat_mxwt[89:72]), (input1_rsci_idat_mxwt[107:90]), (input1_rsci_idat_mxwt[125:108]),
      (input1_rsci_idat_mxwt[143:126]), (input1_rsci_idat_mxwt[161:144]), (input1_rsci_idat_mxwt[179:162]),
      (input1_rsci_idat_mxwt[197:180]), (input1_rsci_idat_mxwt[215:198]), (input1_rsci_idat_mxwt[233:216]),
      (input1_rsci_idat_mxwt[251:234]), (input1_rsci_idat_mxwt[269:252]), (input1_rsci_idat_mxwt[287:270]),
      (input1_rsci_idat_mxwt[305:288]), (input1_rsci_idat_mxwt[323:306]), (input1_rsci_idat_mxwt[341:324]),
      (input1_rsci_idat_mxwt[359:342]), (input1_rsci_idat_mxwt[377:360]), (input1_rsci_idat_mxwt[395:378]),
      (input1_rsci_idat_mxwt[413:396]), (input1_rsci_idat_mxwt[431:414]), (input1_rsci_idat_mxwt[449:432]),
      (input1_rsci_idat_mxwt[467:450]), (input1_rsci_idat_mxwt[485:468]), (input1_rsci_idat_mxwt[503:486]),
      (input1_rsci_idat_mxwt[521:504]), (input1_rsci_idat_mxwt[539:522]), (input1_rsci_idat_mxwt[557:540]),
      (input1_rsci_idat_mxwt[575:558]), (input1_rsci_idat_mxwt[593:576]), (input1_rsci_idat_mxwt[611:594]),
      (input1_rsci_idat_mxwt[629:612]), (input1_rsci_idat_mxwt[647:630]), (input1_rsci_idat_mxwt[665:648]),
      (input1_rsci_idat_mxwt[683:666]), (input1_rsci_idat_mxwt[701:684]), (input1_rsci_idat_mxwt[719:702]),
      (input1_rsci_idat_mxwt[737:720]), (input1_rsci_idat_mxwt[755:738]), (input1_rsci_idat_mxwt[773:756]),
      (input1_rsci_idat_mxwt[791:774]), (input1_rsci_idat_mxwt[809:792]), (input1_rsci_idat_mxwt[827:810]),
      (input1_rsci_idat_mxwt[845:828]), (input1_rsci_idat_mxwt[863:846]), (input1_rsci_idat_mxwt[881:864]),
      (input1_rsci_idat_mxwt[899:882]), (input1_rsci_idat_mxwt[917:900]), (input1_rsci_idat_mxwt[935:918]),
      (input1_rsci_idat_mxwt[953:936]), (input1_rsci_idat_mxwt[971:954]), (input1_rsci_idat_mxwt[989:972]),
      (input1_rsci_idat_mxwt[1007:990]), (input1_rsci_idat_mxwt[1025:1008]), (input1_rsci_idat_mxwt[1043:1026]),
      (input1_rsci_idat_mxwt[1061:1044]), (input1_rsci_idat_mxwt[1079:1062]), (input1_rsci_idat_mxwt[1097:1080]),
      (input1_rsci_idat_mxwt[1115:1098]), (input1_rsci_idat_mxwt[1133:1116]), (input1_rsci_idat_mxwt[1151:1134]),
      (input1_rsci_idat_mxwt[1169:1152]), (input1_rsci_idat_mxwt[1187:1170]), (input1_rsci_idat_mxwt[1205:1188]),
      (input1_rsci_idat_mxwt[1223:1206]), (input1_rsci_idat_mxwt[1241:1224]), (input1_rsci_idat_mxwt[1259:1242]),
      (input1_rsci_idat_mxwt[1277:1260]), (input1_rsci_idat_mxwt[1295:1278]), (input1_rsci_idat_mxwt[1313:1296]),
      (input1_rsci_idat_mxwt[1331:1314]), (input1_rsci_idat_mxwt[1349:1332]), (input1_rsci_idat_mxwt[1367:1350]),
      (input1_rsci_idat_mxwt[1385:1368]), (input1_rsci_idat_mxwt[1403:1386]), (input1_rsci_idat_mxwt[1421:1404]),
      (input1_rsci_idat_mxwt[1439:1422]), (input1_rsci_idat_mxwt[1457:1440]), (input1_rsci_idat_mxwt[1475:1458]),
      (input1_rsci_idat_mxwt[1493:1476]), (input1_rsci_idat_mxwt[1511:1494]), (input1_rsci_idat_mxwt[1529:1512]),
      (input1_rsci_idat_mxwt[1547:1530]), (input1_rsci_idat_mxwt[1565:1548]), (input1_rsci_idat_mxwt[1583:1566]),
      (input1_rsci_idat_mxwt[1601:1584]), (input1_rsci_idat_mxwt[1619:1602]), (input1_rsci_idat_mxwt[1637:1620]),
      (input1_rsci_idat_mxwt[1655:1638]), (input1_rsci_idat_mxwt[1673:1656]), (input1_rsci_idat_mxwt[1691:1674]),
      (input1_rsci_idat_mxwt[1709:1692]), (input1_rsci_idat_mxwt[1727:1710]), (input1_rsci_idat_mxwt[1745:1728]),
      (input1_rsci_idat_mxwt[1763:1746]), (input1_rsci_idat_mxwt[1781:1764]), (input1_rsci_idat_mxwt[1799:1782]),
      (input1_rsci_idat_mxwt[1817:1800]), (input1_rsci_idat_mxwt[1835:1818]), (input1_rsci_idat_mxwt[1853:1836]),
      (input1_rsci_idat_mxwt[1871:1854]), (input1_rsci_idat_mxwt[1889:1872]), (input1_rsci_idat_mxwt[1907:1890]),
      (input1_rsci_idat_mxwt[1925:1908]), (input1_rsci_idat_mxwt[1943:1926]), (input1_rsci_idat_mxwt[1961:1944]),
      (input1_rsci_idat_mxwt[1979:1962]), (input1_rsci_idat_mxwt[1997:1980]), (input1_rsci_idat_mxwt[2015:1998]),
      (input1_rsci_idat_mxwt[2033:2016]), (input1_rsci_idat_mxwt[2051:2034]), (input1_rsci_idat_mxwt[2069:2052]),
      (input1_rsci_idat_mxwt[2087:2070]), (input1_rsci_idat_mxwt[2105:2088]), (input1_rsci_idat_mxwt[2123:2106]),
      (input1_rsci_idat_mxwt[2141:2124]), (input1_rsci_idat_mxwt[2159:2142]), (input1_rsci_idat_mxwt[2177:2160]),
      (input1_rsci_idat_mxwt[2195:2178]), (input1_rsci_idat_mxwt[2213:2196]), (input1_rsci_idat_mxwt[2231:2214]),
      (input1_rsci_idat_mxwt[2249:2232]), (input1_rsci_idat_mxwt[2267:2250]), (input1_rsci_idat_mxwt[2285:2268]),
      (input1_rsci_idat_mxwt[2303:2286]), (input1_rsci_idat_mxwt[2321:2304]), (input1_rsci_idat_mxwt[2339:2322]),
      (input1_rsci_idat_mxwt[2357:2340]), (input1_rsci_idat_mxwt[2375:2358]), (input1_rsci_idat_mxwt[2393:2376]),
      (input1_rsci_idat_mxwt[2411:2394]), (input1_rsci_idat_mxwt[2429:2412]), (input1_rsci_idat_mxwt[2447:2430]),
      (input1_rsci_idat_mxwt[2465:2448]), (input1_rsci_idat_mxwt[2483:2466]), (input1_rsci_idat_mxwt[2501:2484]),
      (input1_rsci_idat_mxwt[2519:2502]), (input1_rsci_idat_mxwt[2537:2520]), (input1_rsci_idat_mxwt[2555:2538]),
      (input1_rsci_idat_mxwt[2573:2556]), (input1_rsci_idat_mxwt[2591:2574]), (input1_rsci_idat_mxwt[2609:2592]),
      (input1_rsci_idat_mxwt[2627:2610]), (input1_rsci_idat_mxwt[2645:2628]), (input1_rsci_idat_mxwt[2663:2646]),
      (input1_rsci_idat_mxwt[2681:2664]), (input1_rsci_idat_mxwt[2699:2682]), (input1_rsci_idat_mxwt[2717:2700]),
      (input1_rsci_idat_mxwt[2735:2718]), (input1_rsci_idat_mxwt[2753:2736]), (input1_rsci_idat_mxwt[2771:2754]),
      (input1_rsci_idat_mxwt[2789:2772]), (input1_rsci_idat_mxwt[2807:2790]), (input1_rsci_idat_mxwt[2825:2808]),
      (input1_rsci_idat_mxwt[2843:2826]), (input1_rsci_idat_mxwt[2861:2844]), (input1_rsci_idat_mxwt[2879:2862]),
      (input1_rsci_idat_mxwt[2897:2880]), (input1_rsci_idat_mxwt[2915:2898]), (input1_rsci_idat_mxwt[2933:2916]),
      (input1_rsci_idat_mxwt[2951:2934]), (input1_rsci_idat_mxwt[2969:2952]), (input1_rsci_idat_mxwt[2987:2970]),
      (input1_rsci_idat_mxwt[3005:2988]), (input1_rsci_idat_mxwt[3023:3006]), (input1_rsci_idat_mxwt[3041:3024]),
      (input1_rsci_idat_mxwt[3059:3042]), (input1_rsci_idat_mxwt[3077:3060]), (input1_rsci_idat_mxwt[3095:3078]),
      (input1_rsci_idat_mxwt[3113:3096]), (input1_rsci_idat_mxwt[3131:3114]), (input1_rsci_idat_mxwt[3149:3132]),
      (input1_rsci_idat_mxwt[3167:3150]), (input1_rsci_idat_mxwt[3185:3168]), (input1_rsci_idat_mxwt[3203:3186]),
      (input1_rsci_idat_mxwt[3221:3204]), (input1_rsci_idat_mxwt[3239:3222]), (input1_rsci_idat_mxwt[3257:3240]),
      (input1_rsci_idat_mxwt[3275:3258]), (input1_rsci_idat_mxwt[3293:3276]), (input1_rsci_idat_mxwt[3311:3294]),
      (input1_rsci_idat_mxwt[3329:3312]), (input1_rsci_idat_mxwt[3347:3330]), (input1_rsci_idat_mxwt[3365:3348]),
      (input1_rsci_idat_mxwt[3383:3366]), (input1_rsci_idat_mxwt[3401:3384]), (input1_rsci_idat_mxwt[3419:3402]),
      (input1_rsci_idat_mxwt[3437:3420]), (input1_rsci_idat_mxwt[3455:3438]), (input1_rsci_idat_mxwt[3473:3456]),
      (input1_rsci_idat_mxwt[3491:3474]), (input1_rsci_idat_mxwt[3509:3492]), (input1_rsci_idat_mxwt[3527:3510]),
      (input1_rsci_idat_mxwt[3545:3528]), (input1_rsci_idat_mxwt[3563:3546]), (input1_rsci_idat_mxwt[3581:3564]),
      (input1_rsci_idat_mxwt[3599:3582]), (input1_rsci_idat_mxwt[3617:3600]), (input1_rsci_idat_mxwt[3635:3618]),
      (input1_rsci_idat_mxwt[3653:3636]), (input1_rsci_idat_mxwt[3671:3654]), (input1_rsci_idat_mxwt[3689:3672]),
      (input1_rsci_idat_mxwt[3707:3690]), (input1_rsci_idat_mxwt[3725:3708]), (input1_rsci_idat_mxwt[3743:3726]),
      (input1_rsci_idat_mxwt[3761:3744]), (input1_rsci_idat_mxwt[3779:3762]), (input1_rsci_idat_mxwt[3797:3780]),
      (input1_rsci_idat_mxwt[3815:3798]), (input1_rsci_idat_mxwt[3833:3816]), (input1_rsci_idat_mxwt[3851:3834]),
      (input1_rsci_idat_mxwt[3869:3852]), (input1_rsci_idat_mxwt[3887:3870]), (input1_rsci_idat_mxwt[3905:3888]),
      (input1_rsci_idat_mxwt[3923:3906]), (input1_rsci_idat_mxwt[3941:3924]), (input1_rsci_idat_mxwt[3959:3942]),
      (input1_rsci_idat_mxwt[3977:3960]), (input1_rsci_idat_mxwt[3995:3978]), (input1_rsci_idat_mxwt[4013:3996]),
      (input1_rsci_idat_mxwt[4031:4014]), (input1_rsci_idat_mxwt[4049:4032]), (input1_rsci_idat_mxwt[4067:4050]),
      (input1_rsci_idat_mxwt[4085:4068]), (input1_rsci_idat_mxwt[4103:4086]), (input1_rsci_idat_mxwt[4121:4104]),
      (input1_rsci_idat_mxwt[4139:4122]), (input1_rsci_idat_mxwt[4157:4140]), (input1_rsci_idat_mxwt[4175:4158]),
      (input1_rsci_idat_mxwt[4193:4176]), (input1_rsci_idat_mxwt[4211:4194]), (input1_rsci_idat_mxwt[4229:4212]),
      (input1_rsci_idat_mxwt[4247:4230]), (input1_rsci_idat_mxwt[4265:4248]), (input1_rsci_idat_mxwt[4283:4266]),
      (input1_rsci_idat_mxwt[4301:4284]), (input1_rsci_idat_mxwt[4319:4302]), (input1_rsci_idat_mxwt[4337:4320]),
      (input1_rsci_idat_mxwt[4355:4338]), (input1_rsci_idat_mxwt[4373:4356]), (input1_rsci_idat_mxwt[4391:4374]),
      (input1_rsci_idat_mxwt[4409:4392]), (input1_rsci_idat_mxwt[4427:4410]), (input1_rsci_idat_mxwt[4445:4428]),
      (input1_rsci_idat_mxwt[4463:4446]), (input1_rsci_idat_mxwt[4481:4464]), (input1_rsci_idat_mxwt[4499:4482]),
      (input1_rsci_idat_mxwt[4517:4500]), (input1_rsci_idat_mxwt[4535:4518]), (input1_rsci_idat_mxwt[4553:4536]),
      (input1_rsci_idat_mxwt[4571:4554]), (input1_rsci_idat_mxwt[4589:4572]), (input1_rsci_idat_mxwt[4607:4590]),
      (input1_rsci_idat_mxwt[4625:4608]), (input1_rsci_idat_mxwt[4643:4626]), (input1_rsci_idat_mxwt[4661:4644]),
      (input1_rsci_idat_mxwt[4679:4662]), (input1_rsci_idat_mxwt[4697:4680]), (input1_rsci_idat_mxwt[4715:4698]),
      (input1_rsci_idat_mxwt[4733:4716]), (input1_rsci_idat_mxwt[4751:4734]), (input1_rsci_idat_mxwt[4769:4752]),
      (input1_rsci_idat_mxwt[4787:4770]), (input1_rsci_idat_mxwt[4805:4788]), (input1_rsci_idat_mxwt[4823:4806]),
      (input1_rsci_idat_mxwt[4841:4824]), (input1_rsci_idat_mxwt[4859:4842]), (input1_rsci_idat_mxwt[4877:4860]),
      (input1_rsci_idat_mxwt[4895:4878]), (input1_rsci_idat_mxwt[4913:4896]), (input1_rsci_idat_mxwt[4931:4914]),
      (input1_rsci_idat_mxwt[4949:4932]), (input1_rsci_idat_mxwt[4967:4950]), (input1_rsci_idat_mxwt[4985:4968]),
      (input1_rsci_idat_mxwt[5003:4986]), (input1_rsci_idat_mxwt[5021:5004]), (input1_rsci_idat_mxwt[5039:5022]),
      (input1_rsci_idat_mxwt[5057:5040]), (input1_rsci_idat_mxwt[5075:5058]), (input1_rsci_idat_mxwt[5093:5076]),
      (input1_rsci_idat_mxwt[5111:5094]), (input1_rsci_idat_mxwt[5129:5112]), (input1_rsci_idat_mxwt[5147:5130]),
      (input1_rsci_idat_mxwt[5165:5148]), (input1_rsci_idat_mxwt[5183:5166]), (input1_rsci_idat_mxwt[5201:5184]),
      (input1_rsci_idat_mxwt[5219:5202]), (input1_rsci_idat_mxwt[5237:5220]), (input1_rsci_idat_mxwt[5255:5238]),
      (input1_rsci_idat_mxwt[5273:5256]), (input1_rsci_idat_mxwt[5291:5274]), (input1_rsci_idat_mxwt[5309:5292]),
      (input1_rsci_idat_mxwt[5327:5310]), (input1_rsci_idat_mxwt[5345:5328]), (input1_rsci_idat_mxwt[5363:5346]),
      (input1_rsci_idat_mxwt[5381:5364]), (input1_rsci_idat_mxwt[5399:5382]), (input1_rsci_idat_mxwt[5417:5400]),
      (input1_rsci_idat_mxwt[5435:5418]), (input1_rsci_idat_mxwt[5453:5436]), (input1_rsci_idat_mxwt[5471:5454]),
      (input1_rsci_idat_mxwt[5489:5472]), (input1_rsci_idat_mxwt[5507:5490]), (input1_rsci_idat_mxwt[5525:5508]),
      (input1_rsci_idat_mxwt[5543:5526]), (input1_rsci_idat_mxwt[5561:5544]), (input1_rsci_idat_mxwt[5579:5562]),
      (input1_rsci_idat_mxwt[5597:5580]), (input1_rsci_idat_mxwt[5615:5598]), (input1_rsci_idat_mxwt[5633:5616]),
      (input1_rsci_idat_mxwt[5651:5634]), (input1_rsci_idat_mxwt[5669:5652]), (input1_rsci_idat_mxwt[5687:5670]),
      (input1_rsci_idat_mxwt[5705:5688]), (input1_rsci_idat_mxwt[5723:5706]), (input1_rsci_idat_mxwt[5741:5724]),
      (input1_rsci_idat_mxwt[5759:5742]), (input1_rsci_idat_mxwt[5777:5760]), (input1_rsci_idat_mxwt[5795:5778]),
      (input1_rsci_idat_mxwt[5813:5796]), (input1_rsci_idat_mxwt[5831:5814]), (input1_rsci_idat_mxwt[5849:5832]),
      (input1_rsci_idat_mxwt[5867:5850]), (input1_rsci_idat_mxwt[5885:5868]), (input1_rsci_idat_mxwt[5903:5886]),
      (input1_rsci_idat_mxwt[5921:5904]), (input1_rsci_idat_mxwt[5939:5922]), (input1_rsci_idat_mxwt[5957:5940]),
      (input1_rsci_idat_mxwt[5975:5958]), (input1_rsci_idat_mxwt[5993:5976]), (input1_rsci_idat_mxwt[6011:5994]),
      (input1_rsci_idat_mxwt[6029:6012]), (input1_rsci_idat_mxwt[6047:6030]), (input1_rsci_idat_mxwt[6065:6048]),
      (input1_rsci_idat_mxwt[6083:6066]), (input1_rsci_idat_mxwt[6101:6084]), (input1_rsci_idat_mxwt[6119:6102]),
      (input1_rsci_idat_mxwt[6137:6120]), (input1_rsci_idat_mxwt[6155:6138]), (input1_rsci_idat_mxwt[6173:6156]),
      (input1_rsci_idat_mxwt[6191:6174]), (input1_rsci_idat_mxwt[6209:6192]), (input1_rsci_idat_mxwt[6227:6210]),
      (input1_rsci_idat_mxwt[6245:6228]), (input1_rsci_idat_mxwt[6263:6246]), (input1_rsci_idat_mxwt[6281:6264]),
      (input1_rsci_idat_mxwt[6299:6282]), (input1_rsci_idat_mxwt[6317:6300]), (input1_rsci_idat_mxwt[6335:6318]),
      (input1_rsci_idat_mxwt[6353:6336]), (input1_rsci_idat_mxwt[6371:6354]), (input1_rsci_idat_mxwt[6389:6372]),
      (input1_rsci_idat_mxwt[6407:6390]), (input1_rsci_idat_mxwt[6425:6408]), (input1_rsci_idat_mxwt[6443:6426]),
      (input1_rsci_idat_mxwt[6461:6444]), (input1_rsci_idat_mxwt[6479:6462]), (input1_rsci_idat_mxwt[6497:6480]),
      (input1_rsci_idat_mxwt[6515:6498]), (input1_rsci_idat_mxwt[6533:6516]), (input1_rsci_idat_mxwt[6551:6534]),
      (input1_rsci_idat_mxwt[6569:6552]), (input1_rsci_idat_mxwt[6587:6570]), (input1_rsci_idat_mxwt[6605:6588]),
      (input1_rsci_idat_mxwt[6623:6606]), (input1_rsci_idat_mxwt[6641:6624]), (input1_rsci_idat_mxwt[6659:6642]),
      (input1_rsci_idat_mxwt[6677:6660]), (input1_rsci_idat_mxwt[6695:6678]), (input1_rsci_idat_mxwt[6713:6696]),
      (input1_rsci_idat_mxwt[6731:6714]), (input1_rsci_idat_mxwt[6749:6732]), (input1_rsci_idat_mxwt[6767:6750]),
      (input1_rsci_idat_mxwt[6785:6768]), (input1_rsci_idat_mxwt[6803:6786]), (input1_rsci_idat_mxwt[6821:6804]),
      (input1_rsci_idat_mxwt[6839:6822]), (input1_rsci_idat_mxwt[6857:6840]), (input1_rsci_idat_mxwt[6875:6858]),
      (input1_rsci_idat_mxwt[6893:6876]), (input1_rsci_idat_mxwt[6911:6894]), (input1_rsci_idat_mxwt[6929:6912]),
      (input1_rsci_idat_mxwt[6947:6930]), (input1_rsci_idat_mxwt[6965:6948]), (input1_rsci_idat_mxwt[6983:6966]),
      (input1_rsci_idat_mxwt[7001:6984]), (input1_rsci_idat_mxwt[7019:7002]), (input1_rsci_idat_mxwt[7037:7020]),
      (input1_rsci_idat_mxwt[7055:7038]), (input1_rsci_idat_mxwt[7073:7056]), (input1_rsci_idat_mxwt[7091:7074]),
      (input1_rsci_idat_mxwt[7109:7092]), (input1_rsci_idat_mxwt[7127:7110]), (input1_rsci_idat_mxwt[7145:7128]),
      (input1_rsci_idat_mxwt[7163:7146]), (input1_rsci_idat_mxwt[7181:7164]), (input1_rsci_idat_mxwt[7199:7182]),
      (input1_rsci_idat_mxwt[7217:7200]), (input1_rsci_idat_mxwt[7235:7218]), (input1_rsci_idat_mxwt[7253:7236]),
      (input1_rsci_idat_mxwt[7271:7254]), (input1_rsci_idat_mxwt[7289:7272]), (input1_rsci_idat_mxwt[7307:7290]),
      (input1_rsci_idat_mxwt[7325:7308]), (input1_rsci_idat_mxwt[7343:7326]), (input1_rsci_idat_mxwt[7361:7344]),
      (input1_rsci_idat_mxwt[7379:7362]), (input1_rsci_idat_mxwt[7397:7380]), (input1_rsci_idat_mxwt[7415:7398]),
      (input1_rsci_idat_mxwt[7433:7416]), (input1_rsci_idat_mxwt[7451:7434]), (input1_rsci_idat_mxwt[7469:7452]),
      (input1_rsci_idat_mxwt[7487:7470]), (input1_rsci_idat_mxwt[7505:7488]), (input1_rsci_idat_mxwt[7523:7506]),
      (input1_rsci_idat_mxwt[7541:7524]), (input1_rsci_idat_mxwt[7559:7542]), (input1_rsci_idat_mxwt[7577:7560]),
      (input1_rsci_idat_mxwt[7595:7578]), (input1_rsci_idat_mxwt[7613:7596]), (input1_rsci_idat_mxwt[7631:7614]),
      (input1_rsci_idat_mxwt[7649:7632]), (input1_rsci_idat_mxwt[7667:7650]), (input1_rsci_idat_mxwt[7685:7668]),
      (input1_rsci_idat_mxwt[7703:7686]), (input1_rsci_idat_mxwt[7721:7704]), (input1_rsci_idat_mxwt[7739:7722]),
      (input1_rsci_idat_mxwt[7757:7740]), (input1_rsci_idat_mxwt[7775:7758]), (input1_rsci_idat_mxwt[7793:7776]),
      (input1_rsci_idat_mxwt[7811:7794]), (input1_rsci_idat_mxwt[7829:7812]), (input1_rsci_idat_mxwt[7847:7830]),
      (input1_rsci_idat_mxwt[7865:7848]), (input1_rsci_idat_mxwt[7883:7866]), (input1_rsci_idat_mxwt[7901:7884]),
      (input1_rsci_idat_mxwt[7919:7902]), (input1_rsci_idat_mxwt[7937:7920]), (input1_rsci_idat_mxwt[7955:7938]),
      (input1_rsci_idat_mxwt[7973:7956]), (input1_rsci_idat_mxwt[7991:7974]), (input1_rsci_idat_mxwt[8009:7992]),
      (input1_rsci_idat_mxwt[8027:8010]), (input1_rsci_idat_mxwt[8045:8028]), (input1_rsci_idat_mxwt[8063:8046]),
      (input1_rsci_idat_mxwt[8081:8064]), (input1_rsci_idat_mxwt[8099:8082]), (input1_rsci_idat_mxwt[8117:8100]),
      (input1_rsci_idat_mxwt[8135:8118]), (input1_rsci_idat_mxwt[8153:8136]), (input1_rsci_idat_mxwt[8171:8154]),
      (input1_rsci_idat_mxwt[8189:8172]), (input1_rsci_idat_mxwt[8207:8190]), (input1_rsci_idat_mxwt[8225:8208]),
      (input1_rsci_idat_mxwt[8243:8226]), (input1_rsci_idat_mxwt[8261:8244]), (input1_rsci_idat_mxwt[8279:8262]),
      (input1_rsci_idat_mxwt[8297:8280]), (input1_rsci_idat_mxwt[8315:8298]), (input1_rsci_idat_mxwt[8333:8316]),
      (input1_rsci_idat_mxwt[8351:8334]), (input1_rsci_idat_mxwt[8369:8352]), (input1_rsci_idat_mxwt[8387:8370]),
      (input1_rsci_idat_mxwt[8405:8388]), (input1_rsci_idat_mxwt[8423:8406]), (input1_rsci_idat_mxwt[8441:8424]),
      (input1_rsci_idat_mxwt[8459:8442]), (input1_rsci_idat_mxwt[8477:8460]), (input1_rsci_idat_mxwt[8495:8478]),
      (input1_rsci_idat_mxwt[8513:8496]), (input1_rsci_idat_mxwt[8531:8514]), (input1_rsci_idat_mxwt[8549:8532]),
      (input1_rsci_idat_mxwt[8567:8550]), (input1_rsci_idat_mxwt[8585:8568]), (input1_rsci_idat_mxwt[8603:8586]),
      (input1_rsci_idat_mxwt[8621:8604]), (input1_rsci_idat_mxwt[8639:8622]), (input1_rsci_idat_mxwt[8657:8640]),
      (input1_rsci_idat_mxwt[8675:8658]), (input1_rsci_idat_mxwt[8693:8676]), (input1_rsci_idat_mxwt[8711:8694]),
      (input1_rsci_idat_mxwt[8729:8712]), (input1_rsci_idat_mxwt[8747:8730]), (input1_rsci_idat_mxwt[8765:8748]),
      (input1_rsci_idat_mxwt[8783:8766]), (input1_rsci_idat_mxwt[8801:8784]), (input1_rsci_idat_mxwt[8819:8802]),
      (input1_rsci_idat_mxwt[8837:8820]), (input1_rsci_idat_mxwt[8855:8838]), (input1_rsci_idat_mxwt[8873:8856]),
      (input1_rsci_idat_mxwt[8891:8874]), (input1_rsci_idat_mxwt[8909:8892]), (input1_rsci_idat_mxwt[8927:8910]),
      (input1_rsci_idat_mxwt[8945:8928]), (input1_rsci_idat_mxwt[8963:8946]), (input1_rsci_idat_mxwt[8981:8964]),
      (input1_rsci_idat_mxwt[8999:8982]), (input1_rsci_idat_mxwt[9017:9000]), (input1_rsci_idat_mxwt[9035:9018]),
      (input1_rsci_idat_mxwt[9053:9036]), (input1_rsci_idat_mxwt[9071:9054]), (input1_rsci_idat_mxwt[9089:9072]),
      (input1_rsci_idat_mxwt[9107:9090]), (input1_rsci_idat_mxwt[9125:9108]), (input1_rsci_idat_mxwt[9143:9126]),
      (input1_rsci_idat_mxwt[9161:9144]), (input1_rsci_idat_mxwt[9179:9162]), (input1_rsci_idat_mxwt[9197:9180]),
      (input1_rsci_idat_mxwt[9215:9198]), (input1_rsci_idat_mxwt[9233:9216]), (input1_rsci_idat_mxwt[9251:9234]),
      (input1_rsci_idat_mxwt[9269:9252]), (input1_rsci_idat_mxwt[9287:9270]), (input1_rsci_idat_mxwt[9305:9288]),
      (input1_rsci_idat_mxwt[9323:9306]), (input1_rsci_idat_mxwt[9341:9324]), (input1_rsci_idat_mxwt[9359:9342]),
      (input1_rsci_idat_mxwt[9377:9360]), (input1_rsci_idat_mxwt[9395:9378]), (input1_rsci_idat_mxwt[9413:9396]),
      (input1_rsci_idat_mxwt[9431:9414]), (input1_rsci_idat_mxwt[9449:9432]), (input1_rsci_idat_mxwt[9467:9450]),
      (input1_rsci_idat_mxwt[9485:9468]), (input1_rsci_idat_mxwt[9503:9486]), (input1_rsci_idat_mxwt[9521:9504]),
      (input1_rsci_idat_mxwt[9539:9522]), (input1_rsci_idat_mxwt[9557:9540]), (input1_rsci_idat_mxwt[9575:9558]),
      (input1_rsci_idat_mxwt[9593:9576]), (input1_rsci_idat_mxwt[9611:9594]), (input1_rsci_idat_mxwt[9629:9612]),
      (input1_rsci_idat_mxwt[9647:9630]), (input1_rsci_idat_mxwt[9665:9648]), (input1_rsci_idat_mxwt[9683:9666]),
      (input1_rsci_idat_mxwt[9701:9684]), (input1_rsci_idat_mxwt[9719:9702]), (input1_rsci_idat_mxwt[9737:9720]),
      (input1_rsci_idat_mxwt[9755:9738]), (input1_rsci_idat_mxwt[9773:9756]), (input1_rsci_idat_mxwt[9791:9774]),
      (input1_rsci_idat_mxwt[9809:9792]), (input1_rsci_idat_mxwt[9827:9810]), (input1_rsci_idat_mxwt[9845:9828]),
      (input1_rsci_idat_mxwt[9863:9846]), (input1_rsci_idat_mxwt[9881:9864]), (input1_rsci_idat_mxwt[9899:9882]),
      (input1_rsci_idat_mxwt[9917:9900]), (input1_rsci_idat_mxwt[9935:9918]), (input1_rsci_idat_mxwt[9953:9936]),
      (input1_rsci_idat_mxwt[9971:9954]), (input1_rsci_idat_mxwt[9989:9972]), (input1_rsci_idat_mxwt[10007:9990]),
      (input1_rsci_idat_mxwt[10025:10008]), (input1_rsci_idat_mxwt[10043:10026]),
      (input1_rsci_idat_mxwt[10061:10044]), (input1_rsci_idat_mxwt[10079:10062]),
      (input1_rsci_idat_mxwt[10097:10080]), (input1_rsci_idat_mxwt[10115:10098]),
      (input1_rsci_idat_mxwt[10133:10116]), (input1_rsci_idat_mxwt[10151:10134]),
      (input1_rsci_idat_mxwt[10169:10152]), (input1_rsci_idat_mxwt[10187:10170]),
      (input1_rsci_idat_mxwt[10205:10188]), (input1_rsci_idat_mxwt[10223:10206]),
      (input1_rsci_idat_mxwt[10241:10224]), (input1_rsci_idat_mxwt[10259:10242]),
      (input1_rsci_idat_mxwt[10277:10260]), (input1_rsci_idat_mxwt[10295:10278]),
      (input1_rsci_idat_mxwt[10313:10296]), (input1_rsci_idat_mxwt[10331:10314]),
      (input1_rsci_idat_mxwt[10349:10332]), (input1_rsci_idat_mxwt[10367:10350]),
      (input1_rsci_idat_mxwt[10385:10368]), (input1_rsci_idat_mxwt[10403:10386]),
      (input1_rsci_idat_mxwt[10421:10404]), (input1_rsci_idat_mxwt[10439:10422]),
      (input1_rsci_idat_mxwt[10457:10440]), (input1_rsci_idat_mxwt[10475:10458]),
      (input1_rsci_idat_mxwt[10493:10476]), (input1_rsci_idat_mxwt[10511:10494]),
      (input1_rsci_idat_mxwt[10529:10512]), (input1_rsci_idat_mxwt[10547:10530]),
      (input1_rsci_idat_mxwt[10565:10548]), (input1_rsci_idat_mxwt[10583:10566]),
      (input1_rsci_idat_mxwt[10601:10584]), (input1_rsci_idat_mxwt[10619:10602]),
      (input1_rsci_idat_mxwt[10637:10620]), (input1_rsci_idat_mxwt[10655:10638]),
      (input1_rsci_idat_mxwt[10673:10656]), (input1_rsci_idat_mxwt[10691:10674]),
      (input1_rsci_idat_mxwt[10709:10692]), (input1_rsci_idat_mxwt[10727:10710]),
      (input1_rsci_idat_mxwt[10745:10728]), (input1_rsci_idat_mxwt[10763:10746]),
      (input1_rsci_idat_mxwt[10781:10764]), (input1_rsci_idat_mxwt[10799:10782]),
      (input1_rsci_idat_mxwt[10817:10800]), (input1_rsci_idat_mxwt[10835:10818]),
      (input1_rsci_idat_mxwt[10853:10836]), (input1_rsci_idat_mxwt[10871:10854]),
      (input1_rsci_idat_mxwt[10889:10872]), (input1_rsci_idat_mxwt[10907:10890]),
      (input1_rsci_idat_mxwt[10925:10908]), (input1_rsci_idat_mxwt[10943:10926]),
      (input1_rsci_idat_mxwt[10961:10944]), (input1_rsci_idat_mxwt[10979:10962]),
      (input1_rsci_idat_mxwt[10997:10980]), (input1_rsci_idat_mxwt[11015:10998]),
      (input1_rsci_idat_mxwt[11033:11016]), (input1_rsci_idat_mxwt[11051:11034]),
      (input1_rsci_idat_mxwt[11069:11052]), (input1_rsci_idat_mxwt[11087:11070]),
      (input1_rsci_idat_mxwt[11105:11088]), (input1_rsci_idat_mxwt[11123:11106]),
      (input1_rsci_idat_mxwt[11141:11124]), (input1_rsci_idat_mxwt[11159:11142]),
      (input1_rsci_idat_mxwt[11177:11160]), (input1_rsci_idat_mxwt[11195:11178]),
      (input1_rsci_idat_mxwt[11213:11196]), (input1_rsci_idat_mxwt[11231:11214]),
      (input1_rsci_idat_mxwt[11249:11232]), (input1_rsci_idat_mxwt[11267:11250]),
      (input1_rsci_idat_mxwt[11285:11268]), (input1_rsci_idat_mxwt[11303:11286]),
      (input1_rsci_idat_mxwt[11321:11304]), (input1_rsci_idat_mxwt[11339:11322]),
      (input1_rsci_idat_mxwt[11357:11340]), (input1_rsci_idat_mxwt[11375:11358]),
      (input1_rsci_idat_mxwt[11393:11376]), (input1_rsci_idat_mxwt[11411:11394]),
      (input1_rsci_idat_mxwt[11429:11412]), (input1_rsci_idat_mxwt[11447:11430]),
      (input1_rsci_idat_mxwt[11465:11448]), (input1_rsci_idat_mxwt[11483:11466]),
      (input1_rsci_idat_mxwt[11501:11484]), (input1_rsci_idat_mxwt[11519:11502]),
      (input1_rsci_idat_mxwt[11537:11520]), (input1_rsci_idat_mxwt[11555:11538]),
      (input1_rsci_idat_mxwt[11573:11556]), (input1_rsci_idat_mxwt[11591:11574]),
      (input1_rsci_idat_mxwt[11609:11592]), (input1_rsci_idat_mxwt[11627:11610]),
      (input1_rsci_idat_mxwt[11645:11628]), (input1_rsci_idat_mxwt[11663:11646]),
      (input1_rsci_idat_mxwt[11681:11664]), (input1_rsci_idat_mxwt[11699:11682]),
      (input1_rsci_idat_mxwt[11717:11700]), (input1_rsci_idat_mxwt[11735:11718]),
      (input1_rsci_idat_mxwt[11753:11736]), (input1_rsci_idat_mxwt[11771:11754]),
      (input1_rsci_idat_mxwt[11789:11772]), (input1_rsci_idat_mxwt[11807:11790]),
      (input1_rsci_idat_mxwt[11825:11808]), (input1_rsci_idat_mxwt[11843:11826]),
      (input1_rsci_idat_mxwt[11861:11844]), (input1_rsci_idat_mxwt[11879:11862]),
      (input1_rsci_idat_mxwt[11897:11880]), (input1_rsci_idat_mxwt[11915:11898]),
      (input1_rsci_idat_mxwt[11933:11916]), (input1_rsci_idat_mxwt[11951:11934]),
      (input1_rsci_idat_mxwt[11969:11952]), (input1_rsci_idat_mxwt[11987:11970]),
      (input1_rsci_idat_mxwt[12005:11988]), (input1_rsci_idat_mxwt[12023:12006]),
      (input1_rsci_idat_mxwt[12041:12024]), (input1_rsci_idat_mxwt[12059:12042]),
      (input1_rsci_idat_mxwt[12077:12060]), (input1_rsci_idat_mxwt[12095:12078]),
      (input1_rsci_idat_mxwt[12113:12096]), (input1_rsci_idat_mxwt[12131:12114]),
      (input1_rsci_idat_mxwt[12149:12132]), (input1_rsci_idat_mxwt[12167:12150]),
      (input1_rsci_idat_mxwt[12185:12168]), (input1_rsci_idat_mxwt[12203:12186]),
      (input1_rsci_idat_mxwt[12221:12204]), (input1_rsci_idat_mxwt[12239:12222]),
      (input1_rsci_idat_mxwt[12257:12240]), (input1_rsci_idat_mxwt[12275:12258]),
      (input1_rsci_idat_mxwt[12293:12276]), (input1_rsci_idat_mxwt[12311:12294]),
      (input1_rsci_idat_mxwt[12329:12312]), (input1_rsci_idat_mxwt[12347:12330]),
      (input1_rsci_idat_mxwt[12365:12348]), (input1_rsci_idat_mxwt[12383:12366]),
      (input1_rsci_idat_mxwt[12401:12384]), (input1_rsci_idat_mxwt[12419:12402]),
      (input1_rsci_idat_mxwt[12437:12420]), (input1_rsci_idat_mxwt[12455:12438]),
      (input1_rsci_idat_mxwt[12473:12456]), (input1_rsci_idat_mxwt[12491:12474]),
      (input1_rsci_idat_mxwt[12509:12492]), (input1_rsci_idat_mxwt[12527:12510]),
      (input1_rsci_idat_mxwt[12545:12528]), (input1_rsci_idat_mxwt[12563:12546]),
      (input1_rsci_idat_mxwt[12581:12564]), (input1_rsci_idat_mxwt[12599:12582]),
      (input1_rsci_idat_mxwt[12617:12600]), (input1_rsci_idat_mxwt[12635:12618]),
      (input1_rsci_idat_mxwt[12653:12636]), (input1_rsci_idat_mxwt[12671:12654]),
      (input1_rsci_idat_mxwt[12689:12672]), (input1_rsci_idat_mxwt[12707:12690]),
      (input1_rsci_idat_mxwt[12725:12708]), (input1_rsci_idat_mxwt[12743:12726]),
      (input1_rsci_idat_mxwt[12761:12744]), (input1_rsci_idat_mxwt[12779:12762]),
      (input1_rsci_idat_mxwt[12797:12780]), (input1_rsci_idat_mxwt[12815:12798]),
      (input1_rsci_idat_mxwt[12833:12816]), (input1_rsci_idat_mxwt[12851:12834]),
      (input1_rsci_idat_mxwt[12869:12852]), (input1_rsci_idat_mxwt[12887:12870]),
      (input1_rsci_idat_mxwt[12905:12888]), (input1_rsci_idat_mxwt[12923:12906]),
      (input1_rsci_idat_mxwt[12941:12924]), (input1_rsci_idat_mxwt[12959:12942]),
      (input1_rsci_idat_mxwt[12977:12960]), (input1_rsci_idat_mxwt[12995:12978]),
      (input1_rsci_idat_mxwt[13013:12996]), (input1_rsci_idat_mxwt[13031:13014]),
      (input1_rsci_idat_mxwt[13049:13032]), (input1_rsci_idat_mxwt[13067:13050]),
      (input1_rsci_idat_mxwt[13085:13068]), (input1_rsci_idat_mxwt[13103:13086]),
      (input1_rsci_idat_mxwt[13121:13104]), (input1_rsci_idat_mxwt[13139:13122]),
      (input1_rsci_idat_mxwt[13157:13140]), (input1_rsci_idat_mxwt[13175:13158]),
      (input1_rsci_idat_mxwt[13193:13176]), (input1_rsci_idat_mxwt[13211:13194]),
      (input1_rsci_idat_mxwt[13229:13212]), (input1_rsci_idat_mxwt[13247:13230]),
      (input1_rsci_idat_mxwt[13265:13248]), (input1_rsci_idat_mxwt[13283:13266]),
      (input1_rsci_idat_mxwt[13301:13284]), (input1_rsci_idat_mxwt[13319:13302]),
      (input1_rsci_idat_mxwt[13337:13320]), (input1_rsci_idat_mxwt[13355:13338]),
      (input1_rsci_idat_mxwt[13373:13356]), (input1_rsci_idat_mxwt[13391:13374]),
      (input1_rsci_idat_mxwt[13409:13392]), (input1_rsci_idat_mxwt[13427:13410]),
      (input1_rsci_idat_mxwt[13445:13428]), (input1_rsci_idat_mxwt[13463:13446]),
      (input1_rsci_idat_mxwt[13481:13464]), (input1_rsci_idat_mxwt[13499:13482]),
      (input1_rsci_idat_mxwt[13517:13500]), (input1_rsci_idat_mxwt[13535:13518]),
      (input1_rsci_idat_mxwt[13553:13536]), (input1_rsci_idat_mxwt[13571:13554]),
      (input1_rsci_idat_mxwt[13589:13572]), (input1_rsci_idat_mxwt[13607:13590]),
      (input1_rsci_idat_mxwt[13625:13608]), (input1_rsci_idat_mxwt[13643:13626]),
      (input1_rsci_idat_mxwt[13661:13644]), (input1_rsci_idat_mxwt[13679:13662]),
      (input1_rsci_idat_mxwt[13697:13680]), (input1_rsci_idat_mxwt[13715:13698]),
      (input1_rsci_idat_mxwt[13733:13716]), (input1_rsci_idat_mxwt[13751:13734]),
      (input1_rsci_idat_mxwt[13769:13752]), (input1_rsci_idat_mxwt[13787:13770]),
      (input1_rsci_idat_mxwt[13805:13788]), (input1_rsci_idat_mxwt[13823:13806]),
      (input1_rsci_idat_mxwt[13841:13824]), (input1_rsci_idat_mxwt[13859:13842]),
      (input1_rsci_idat_mxwt[13877:13860]), (input1_rsci_idat_mxwt[13895:13878]),
      (input1_rsci_idat_mxwt[13913:13896]), (input1_rsci_idat_mxwt[13931:13914]),
      (input1_rsci_idat_mxwt[13949:13932]), (input1_rsci_idat_mxwt[13967:13950]),
      (input1_rsci_idat_mxwt[13985:13968]), (input1_rsci_idat_mxwt[14003:13986]),
      (input1_rsci_idat_mxwt[14021:14004]), (input1_rsci_idat_mxwt[14039:14022]),
      (input1_rsci_idat_mxwt[14057:14040]), (input1_rsci_idat_mxwt[14075:14058]),
      (input1_rsci_idat_mxwt[14093:14076]), (input1_rsci_idat_mxwt[14111:14094]),
      layer3_out_0_16_0_lpi_1_dfm_11_0[9:0]);
  assign nl_IndexLoop_if_acc_13_nl = conv_u2s_5_6({(IndexLoop_if_acc_3_psp_1_sva_1[7])
      , 1'b0 , (signext_2_1(IndexLoop_if_acc_3_psp_1_sva_1[7])) , 1'b1}) + conv_u2s_5_6({4'b1110
      , (~ (IndexLoop_if_acc_3_psp_1_sva_1[6]))});
  assign IndexLoop_if_acc_13_nl = nl_IndexLoop_if_acc_13_nl[5:0];
  assign nl_IndexLoop_if_acc_15_nl = ({1'b1 , (~ (IndexLoop_if_acc_3_psp_1_sva_1[5]))})
      + 2'b11;
  assign IndexLoop_if_acc_15_nl = nl_IndexLoop_if_acc_15_nl[1:0];
  assign nl_IndexLoop_if_acc_10_nl = conv_u2u_6_7({(z_out[1:0]) , (IndexLoop_if_acc_3_psp_1_sva_1[7])
      , (IndexLoop_if_acc_3_psp_1_sva_1[7]) , (IndexLoop_if_acc_15_nl)}) + conv_u2u_5_7(IndexLoop_if_acc_3_psp_1_sva_1[4:0]);
  assign IndexLoop_if_acc_10_nl = nl_IndexLoop_if_acc_10_nl[6:0];
  assign nl_IndexLoop_if_acc_4_psp_sva_1 = ({(~ (IndexLoop_if_acc_3_psp_1_sva_1[7]))
      , (IndexLoop_if_acc_13_nl)}) + (IndexLoop_if_acc_10_nl);
  assign IndexLoop_if_acc_4_psp_sva_1 = nl_IndexLoop_if_acc_4_psp_sva_1[6:0];
  assign nl_IndexLoop_if_acc_12_nl = conv_u2u_3_4({(z_out_13[10]) , (signext_2_1(z_out_13[11]))})
      + conv_u2u_1_4(~ (z_out_13[14])) + 4'b0001;
  assign IndexLoop_if_acc_12_nl = nl_IndexLoop_if_acc_12_nl[3:0];
  assign nl_IndexLoop_if_acc_8_nl = conv_u2u_6_8({(IndexLoop_if_acc_12_nl) , (~ (z_out_13[13:12]))})
      + conv_u2u_6_8({(z_out_13[13:12]) , 3'b000 , (z_out_13[11])}) + conv_u2u_6_8({(~
      (z_out_13[11])) , (~ (z_out_13[9])) , (~ (z_out_13[13:12])) , 1'b1 , (~ (z_out_13[9]))})
      + conv_u2u_5_8(z_out_13[8:4]) + conv_u2u_1_8(~ (z_out_13[14]));
  assign IndexLoop_if_acc_8_nl = nl_IndexLoop_if_acc_8_nl[7:0];
  assign nl_IndexLoop_if_acc_3_psp_1_sva_1 = (IndexLoop_if_acc_8_nl) + ({7'b1011010
      , (~ (z_out_13[10]))});
  assign IndexLoop_if_acc_3_psp_1_sva_1 = nl_IndexLoop_if_acc_3_psp_1_sva_1[7:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_63_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_16_0_lpi_1_dfm_mx0w2
      = MUX_v_17_2_2(17'b00000000000000000, (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_63_sva[16:0]),
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_16_0_lpi_1_dfm_mx0w2
      = MUX_v_17_2_2(17'b00000000000000000, (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_61_1_sva_2[16:0]),
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12
      = MUX_v_5_2_2(5'b00000, (reg_MultLoop_1_mux_64_itm_1_reg[4:0]), (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0
      = MUX_v_12_2_2(12'b000000000000, reg_MultLoop_1_mux_64_itm_1_1_reg, (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
      = MUX_v_2_2_2(2'b00, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_16_15,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0
      = MUX_v_15_2_2(15'b000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_14_0,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_16_0_lpi_1_dfm_mx0w2_16_15
      = MUX_v_2_2_2(2'b00, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_16_15,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_16_0_lpi_1_dfm_mx0w2_14_0
      = MUX_v_15_2_2(15'b000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_14_0,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_16_0_lpi_1_dfm_mx0w2
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_16_0_lpi_1_dfm_mx0w2
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_16_0_lpi_1_dfm_mx0w2
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_6_1_sva_2[16:0]),
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_16_0_lpi_1_dfm_mx0w2
      = MUX_v_17_2_2(17'b00000000000000000, (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_59_1_sva_2[16:0]),
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12
      = MUX_v_5_2_2(5'b00000, (reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_reg[4:0]),
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0
      = MUX_v_12_2_2(12'b000000000000, reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_1_reg,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12
      = MUX_v_5_2_2(5'b00000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_2_reg,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_10
      = MUX_v_2_2_2(2'b00, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_4_reg,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_9_0
      = MUX_v_10_2_2(10'b0000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd_2,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12
      = MUX_v_5_2_2(5'b00000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_2_reg,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0
      = MUX_v_12_2_2(12'b000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_3_reg,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12
      = MUX_v_5_2_2(5'b00000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_2_reg,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0
      = MUX_v_12_2_2(12'b000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_3_reg,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12
      = MUX_v_5_2_2(5'b00000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_2_reg,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0
      = MUX_v_12_2_2(12'b000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_3_reg,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2[16:0]),
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
      = MUX_v_2_2_2(2'b00, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_16_15,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0
      = MUX_v_15_2_2(15'b000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_14_0,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
      = MUX_v_2_2_2(2'b00, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_16_15,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0
      = MUX_v_15_2_2(15'b000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_14_0,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
      = MUX_v_2_2_2(2'b00, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_16_15,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0
      = MUX_v_15_2_2(15'b000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_14_0,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
      = MUX_v_2_2_2(2'b00, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_16_15,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0
      = MUX_v_15_2_2(15'b000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_14_0,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
      = MUX_v_2_2_2(2'b00, (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_1_ftd[1:0]),
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_12
      = MUX_v_3_2_2(3'b000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_2_reg,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0
      = MUX_v_12_2_2(12'b000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
      = MUX_v_2_2_2(2'b00, (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd[1:0]),
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_12
      = MUX_v_3_2_2(3'b000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_2_reg,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11
      = reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_4_reg
      & (z_out_23_22_8[10]);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_10_0
      = MUX_v_11_2_2(11'b00000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_1_ftd_1,
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_58_1_sva_2[16:0]),
      (z_out_23_22_8[10]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_16_0_lpi_1_dfm_mx0w0
      = MUX_v_17_2_2(17'b00000000000000000, (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_60_1_sva_2[16:0]),
      (z_out_23_22_8[10]));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_4_sva_mx0w1
      = ~(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd
      | (~((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_2_reg[4:3]!=2'b00))));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_3_sva_mx0w1
      = ~((reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_reg[5])
      | (~((reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_reg[4:3]!=2'b00))));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_2_sva_mx0w1
      = ~((reg_MultLoop_1_mux_64_itm_1_reg[5]) | (~((reg_MultLoop_1_mux_64_itm_1_reg[4:3]!=2'b00))));
  assign nl_MultLoop_2_1_acc_3_tmp = ROM_1i9_1o3_2fa806bf16b3e0d54016201674d036b62f_1
      + 3'b101;
  assign MultLoop_2_1_acc_3_tmp = nl_MultLoop_2_1_acc_3_tmp[2:0];
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_sva_mx0w0 =
      ~((nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2[17])
      | (~((nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2[16:15]!=2'b00))));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_9_sva_mx0w0
      = ~(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd
      | (~((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd_1[16:15]!=2'b00))));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_8_sva_mx0w0
      = ~(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd
      | (~((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd_1[16:15]!=2'b00))));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_7_sva_mx0w0
      = ~(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_1_ftd
      | (~((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_2_reg[4:3]!=2'b00))));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_6_sva_mx0w0
      = ~(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_1_ftd
      | (~((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_2_reg[4:3]!=2'b00))));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_5_sva_mx0w0
      = ~(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_1_ftd
      | (~((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_2_reg[4:3]!=2'b00))));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_1_nor_2_nl = ~(MUX_v_15_2_2(({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_1_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_2_reg}),
      15'b111111111111111, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_1_sva_1));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_1_and_nl = (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg[2])
      & (~((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg[1:0]==2'b11)));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_1_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_psp_sva_1
      = ~(MUX_v_15_2_2((nnet_softmax_layer6_t_result_t_softmax_config7_for_1_nor_2_nl),
      15'b111111111111111, (nnet_softmax_layer6_t_result_t_softmax_config7_for_1_and_nl)));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_1_sva_1 = ~((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg[2])
      | (~((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg[1:0]!=2'b00))));
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000
      = MUX_v_12_10_2(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg,
      reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_1_reg,
      reg_MultLoop_1_mux_64_itm_1_1_reg, layer3_out_0_16_0_lpi_1_dfm_11_0, ({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_4_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2}),
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_2_reg,
      ({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_4_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd_2}),
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_3_reg,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_3_reg,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_3_reg,
      InitAccumLoop_2_iacc_3_0_sva);
  assign nnet_softmax_layer6_t_result_t_softmax_config7_for_1_or_tmp = (InitAccumLoop_2_iacc_3_0_sva!=4'b0000);
  assign and_dcpl = ~((fsm_output[6:5]!=2'b00));
  assign or_tmp_1 = (~ (fsm_output[3])) | (fsm_output[4]) | (~ (fsm_output[7]));
  assign or_tmp_2 = (fsm_output[4]) | (~ (fsm_output[7]));
  assign mux_tmp_2 = MUX_s_1_2_2((~ and_2631_cse), or_tmp_2, fsm_output[3]);
  assign mux_33_cse = MUX_s_1_2_2(mux_661_cse, or_864_cse, fsm_output[2]);
  assign or_tmp_48 = nor_943_cse | (fsm_output[7]);
  assign or_1409_nl = (fsm_output[6:4]!=3'b000);
  assign mux_tmp_81 = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), or_1409_nl);
  assign or_tmp_91 = (fsm_output[7:6]!=2'b00);
  assign mux_tmp_183 = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), or_1398_cse);
  assign mux_tmp_184 = MUX_s_1_2_2(mux_tmp_183, or_1213_cse, or_941_cse);
  assign or_tmp_196 = (fsm_output[5]) | mux_661_cse;
  assign or_tmp_231 = (~ (fsm_output[4])) | (~ (fsm_output[5])) | (fsm_output[7]);
  assign or_609_nl = (fsm_output[5:4]!=2'b00) | mux_661_cse;
  assign mux_tmp_377 = MUX_s_1_2_2((or_609_nl), or_tmp_231, fsm_output[3]);
  assign nand_tmp_14 = ~((fsm_output[2]) & (~ mux_661_cse));
  assign mux_tmp_419 = MUX_s_1_2_2(nand_tmp_14, mux_33_cse, fsm_output[1]);
  assign mux_421_cse = MUX_s_1_2_2(or_1298_cse, mux_33_cse, fsm_output[1]);
  assign mux_456_cse = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), fsm_output[2]);
  assign nor_310_cse = ~(and_817_cse | (fsm_output[3]));
  assign and_dcpl_50 = (fsm_output[3:2]==2'b01);
  assign and_dcpl_51 = and_dcpl_50 & and_810_cse_1;
  assign and_dcpl_53 = (fsm_output[7:6]==2'b10);
  assign and_dcpl_54 = and_dcpl_53 & nor_943_cse;
  assign and_dcpl_55 = and_dcpl_54 & and_dcpl_51;
  assign and_dcpl_56 = (fsm_output[1:0]==2'b01);
  assign and_dcpl_57 = and_dcpl_50 & and_dcpl_56;
  assign and_dcpl_58 = (fsm_output[7:6]==2'b01);
  assign and_dcpl_59 = and_dcpl_58 & nor_943_cse;
  assign and_dcpl_60 = and_dcpl_59 & and_dcpl_57;
  assign and_dcpl_62 = nor_942_cse & and_810_cse_1;
  assign and_dcpl_64 = nor_944_cse & nor_943_cse;
  assign and_dcpl_65 = and_dcpl_64 & and_dcpl_62;
  assign and_dcpl_66 = (fsm_output[0]) & IndexLoop_stage_0;
  assign and_dcpl_70 = and_dcpl_53 & (~ (fsm_output[5]));
  assign and_dcpl_73 = (fsm_output[2:1]==2'b10);
  assign and_dcpl_75 = and_dcpl_58 & (~ (fsm_output[5]));
  assign and_dcpl_77 = and_dcpl_75 & nor_298_cse & and_dcpl_73 & and_dcpl_66;
  assign and_dcpl_82 = nor_944_cse & (~ (fsm_output[5])) & nor_298_cse & (fsm_output[2:1]==2'b01)
      & and_dcpl_66;
  assign and_dcpl_84 = and_817_cse & (~ (fsm_output[0]));
  assign and_dcpl_87 = and_dcpl_70 & and_862_cse;
  assign or_dcpl_334 = or_864_cse | (fsm_output[5]);
  assign and_dcpl_92 = ~((InitAccumLoop_2_iacc_3_0_sva[2:1]!=2'b00));
  assign and_dcpl_93 = and_dcpl_92 & (InitAccumLoop_2_iacc_3_0_sva[0]);
  assign and_dcpl_94 = (~ (fsm_output[0])) & IndexLoop_stage_0;
  assign and_dcpl_95 = and_dcpl_94 & (~ (InitAccumLoop_2_iacc_3_0_sva[3]));
  assign and_dcpl_99 = (fsm_output[5:4]==2'b01);
  assign and_dcpl_100 = and_dcpl_53 & and_dcpl_99;
  assign and_dcpl_101 = and_dcpl_100 & and_2650_cse & (fsm_output[1]);
  assign and_dcpl_103 = (fsm_output[1:0]==2'b10);
  assign and_dcpl_106 = and_862_cse & (fsm_output[2]) & and_dcpl_103 & IndexLoop_stage_0;
  assign or_dcpl_337 = (InitAccumLoop_2_iacc_3_0_sva[1:0]!=2'b01);
  assign or_dcpl_338 = (InitAccumLoop_2_iacc_3_0_sva[3:2]!=2'b00);
  assign or_dcpl_339 = or_dcpl_338 | or_dcpl_337;
  assign and_dcpl_109 = (InitAccumLoop_2_iacc_3_0_sva[2:1]==2'b01);
  assign or_dcpl_340 = (InitAccumLoop_2_iacc_3_0_sva[1:0]!=2'b10);
  assign or_dcpl_341 = or_dcpl_338 | or_dcpl_340;
  assign or_dcpl_342 = ~((InitAccumLoop_2_iacc_3_0_sva[1:0]==2'b11));
  assign or_dcpl_343 = or_dcpl_338 | or_dcpl_342;
  assign and_dcpl_120 = (InitAccumLoop_2_iacc_3_0_sva[2:1]==2'b10);
  assign or_dcpl_344 = (InitAccumLoop_2_iacc_3_0_sva[1:0]!=2'b00);
  assign or_dcpl_345 = (InitAccumLoop_2_iacc_3_0_sva[3:2]!=2'b01);
  assign or_dcpl_346 = or_dcpl_345 | or_dcpl_344;
  assign or_dcpl_347 = or_dcpl_345 | or_dcpl_337;
  assign and_dcpl_131 = (InitAccumLoop_2_iacc_3_0_sva[2:1]==2'b11);
  assign or_dcpl_348 = or_dcpl_345 | or_dcpl_340;
  assign or_dcpl_349 = or_dcpl_345 | or_dcpl_342;
  assign and_dcpl_143 = and_dcpl_94 & (InitAccumLoop_2_iacc_3_0_sva[3]);
  assign or_dcpl_350 = (InitAccumLoop_2_iacc_3_0_sva[3:2]!=2'b10);
  assign or_dcpl_351 = or_dcpl_350 | or_dcpl_344;
  assign and_dcpl_154 = nor_942_cse & and_dcpl_103;
  assign and_dcpl_155 = and_dcpl_64 & and_dcpl_154;
  assign or_dcpl_362 = ~((InitAccumLoop_1_iacc_6_0_sva_5_0[2:1]==2'b11));
  assign or_dcpl_363 = or_dcpl_362 | (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[5]));
  assign or_dcpl_364 = (InitAccumLoop_1_iacc_6_0_sva_5_0[0]) | (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[4]));
  assign or_dcpl_365 = or_dcpl_364 | (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[3]));
  assign or_dcpl_366 = or_dcpl_365 | or_dcpl_363;
  assign or_dcpl_368 = (InitAccumLoop_1_iacc_6_0_sva_5_0[2:1]!=2'b00);
  assign or_dcpl_369 = or_dcpl_368 | (InitAccumLoop_1_iacc_6_0_sva_5_0[5]);
  assign or_dcpl_370 = (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[0])) | (InitAccumLoop_1_iacc_6_0_sva_5_0[4]);
  assign or_dcpl_371 = or_dcpl_370 | (InitAccumLoop_1_iacc_6_0_sva_5_0[3]);
  assign or_dcpl_372 = or_dcpl_371 | or_dcpl_369;
  assign or_dcpl_373 = (InitAccumLoop_1_iacc_6_0_sva_5_0[2:1]!=2'b10);
  assign or_dcpl_374 = or_dcpl_373 | (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[5]));
  assign or_dcpl_375 = ~((InitAccumLoop_1_iacc_6_0_sva_5_0[0]) & (InitAccumLoop_1_iacc_6_0_sva_5_0[4]));
  assign or_dcpl_376 = or_dcpl_375 | (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[3]));
  assign or_dcpl_377 = or_dcpl_376 | or_dcpl_374;
  assign or_dcpl_378 = (InitAccumLoop_1_iacc_6_0_sva_5_0[2:1]!=2'b01);
  assign or_dcpl_379 = or_dcpl_378 | (InitAccumLoop_1_iacc_6_0_sva_5_0[5]);
  assign or_dcpl_380 = (InitAccumLoop_1_iacc_6_0_sva_5_0[0]) | (InitAccumLoop_1_iacc_6_0_sva_5_0[4]);
  assign or_dcpl_381 = or_dcpl_380 | (InitAccumLoop_1_iacc_6_0_sva_5_0[3]);
  assign or_dcpl_382 = or_dcpl_381 | or_dcpl_379;
  assign or_dcpl_383 = or_dcpl_365 | or_dcpl_374;
  assign or_dcpl_384 = or_dcpl_371 | or_dcpl_379;
  assign or_dcpl_385 = or_dcpl_378 | (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[5]));
  assign or_dcpl_386 = or_dcpl_376 | or_dcpl_385;
  assign or_dcpl_387 = or_dcpl_373 | (InitAccumLoop_1_iacc_6_0_sva_5_0[5]);
  assign or_dcpl_388 = or_dcpl_381 | or_dcpl_387;
  assign or_dcpl_389 = or_dcpl_365 | or_dcpl_385;
  assign or_dcpl_390 = or_dcpl_371 | or_dcpl_387;
  assign or_dcpl_391 = or_dcpl_368 | (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[5]));
  assign or_dcpl_392 = or_dcpl_376 | or_dcpl_391;
  assign or_dcpl_393 = or_dcpl_362 | (InitAccumLoop_1_iacc_6_0_sva_5_0[5]);
  assign or_dcpl_394 = or_dcpl_381 | or_dcpl_393;
  assign or_dcpl_395 = or_dcpl_365 | or_dcpl_391;
  assign or_dcpl_396 = or_dcpl_371 | or_dcpl_393;
  assign or_dcpl_397 = or_dcpl_375 | (InitAccumLoop_1_iacc_6_0_sva_5_0[3]);
  assign or_dcpl_398 = or_dcpl_397 | or_dcpl_363;
  assign or_dcpl_399 = or_dcpl_380 | (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[3]));
  assign or_dcpl_400 = or_dcpl_399 | or_dcpl_369;
  assign or_dcpl_401 = or_dcpl_364 | (InitAccumLoop_1_iacc_6_0_sva_5_0[3]);
  assign or_dcpl_402 = or_dcpl_401 | or_dcpl_363;
  assign or_dcpl_403 = or_dcpl_370 | (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[3]));
  assign or_dcpl_404 = or_dcpl_403 | or_dcpl_369;
  assign or_dcpl_405 = or_dcpl_397 | or_dcpl_374;
  assign or_dcpl_406 = or_dcpl_399 | or_dcpl_379;
  assign or_dcpl_407 = or_dcpl_401 | or_dcpl_374;
  assign or_dcpl_408 = or_dcpl_403 | or_dcpl_379;
  assign or_dcpl_409 = or_dcpl_397 | or_dcpl_385;
  assign or_dcpl_410 = or_dcpl_399 | or_dcpl_387;
  assign or_dcpl_411 = or_dcpl_401 | or_dcpl_385;
  assign or_dcpl_412 = or_dcpl_403 | or_dcpl_387;
  assign or_dcpl_413 = or_dcpl_397 | or_dcpl_391;
  assign or_dcpl_414 = or_dcpl_399 | or_dcpl_393;
  assign or_dcpl_415 = or_dcpl_401 | or_dcpl_391;
  assign or_dcpl_416 = or_dcpl_403 | or_dcpl_393;
  assign or_dcpl_417 = or_dcpl_403 | or_dcpl_363;
  assign or_dcpl_418 = or_dcpl_401 | or_dcpl_369;
  assign or_dcpl_419 = or_dcpl_399 | or_dcpl_363;
  assign or_dcpl_420 = or_dcpl_397 | or_dcpl_369;
  assign or_dcpl_421 = or_dcpl_403 | or_dcpl_374;
  assign or_dcpl_422 = or_dcpl_401 | or_dcpl_379;
  assign or_dcpl_423 = or_dcpl_399 | or_dcpl_374;
  assign or_dcpl_424 = or_dcpl_397 | or_dcpl_379;
  assign or_dcpl_425 = or_dcpl_403 | or_dcpl_385;
  assign or_dcpl_426 = or_dcpl_401 | or_dcpl_387;
  assign or_dcpl_427 = or_dcpl_399 | or_dcpl_385;
  assign or_dcpl_428 = or_dcpl_397 | or_dcpl_387;
  assign or_dcpl_429 = or_dcpl_403 | or_dcpl_391;
  assign or_dcpl_430 = or_dcpl_401 | or_dcpl_393;
  assign or_dcpl_431 = or_dcpl_399 | or_dcpl_391;
  assign or_dcpl_432 = or_dcpl_397 | or_dcpl_393;
  assign or_dcpl_433 = or_dcpl_371 | or_dcpl_363;
  assign or_dcpl_434 = or_dcpl_365 | or_dcpl_369;
  assign or_dcpl_435 = or_dcpl_381 | or_dcpl_363;
  assign or_dcpl_436 = or_dcpl_376 | or_dcpl_369;
  assign or_dcpl_437 = or_dcpl_371 | or_dcpl_374;
  assign or_dcpl_438 = or_dcpl_365 | or_dcpl_379;
  assign or_dcpl_439 = or_dcpl_381 | or_dcpl_374;
  assign or_dcpl_440 = or_dcpl_376 | or_dcpl_379;
  assign or_dcpl_441 = or_dcpl_371 | or_dcpl_385;
  assign or_dcpl_442 = or_dcpl_365 | or_dcpl_387;
  assign or_dcpl_443 = or_dcpl_381 | or_dcpl_385;
  assign or_dcpl_444 = or_dcpl_376 | or_dcpl_387;
  assign or_dcpl_445 = or_dcpl_371 | or_dcpl_391;
  assign or_dcpl_446 = or_dcpl_365 | or_dcpl_393;
  assign or_dcpl_447 = or_dcpl_381 | or_dcpl_391;
  assign or_dcpl_448 = or_dcpl_376 | or_dcpl_393;
  assign and_dcpl_157 = and_dcpl_50 & nor_306_cse;
  assign and_dcpl_158 = and_dcpl_59 & and_dcpl_157;
  assign and_dcpl_159 = and_dcpl_50 & and_dcpl_103;
  assign and_dcpl_160 = and_dcpl_54 & and_dcpl_159;
  assign or_dcpl_455 = or_864_cse | or_888_cse;
  assign or_dcpl_465 = (fsm_output[1:0]!=2'b10);
  assign or_dcpl_466 = ~((fsm_output[3:2]==2'b11));
  assign or_dcpl_467 = or_dcpl_466 | or_dcpl_465;
  assign or_dcpl_469 = or_864_cse | (fsm_output[5:4]!=2'b01);
  assign or_dcpl_471 = (~ IndexLoop_stage_0) | (InitAccumLoop_2_iacc_3_0_sva[3]);
  assign or_dcpl_472 = or_dcpl_471 | (~ (InitAccumLoop_2_iacc_3_0_sva[2]));
  assign or_dcpl_481 = (~ IndexLoop_stage_0) | (InitAccumLoop_2_iacc_3_0_sva[3:2]!=2'b10);
  assign or_dcpl_484 = or_dcpl_471 | (InitAccumLoop_2_iacc_3_0_sva[2]);
  assign and_dcpl_169 = nor_943_cse & (~ (fsm_output[3]));
  assign and_dcpl_171 = (fsm_output[3:2]==2'b10);
  assign mux_479_nl = MUX_s_1_2_2(or_10_cse, (~ and_817_cse), fsm_output[0]);
  assign and_dcpl_175 = and_dcpl_100 & (mux_479_nl) & (fsm_output[3]);
  assign or_dcpl_490 = or_dcpl_381 | or_dcpl_369;
  assign and_dcpl_176 = (~ IndexLoop_stage_0) & IndexLoop_stage_0_2;
  assign and_dcpl_177 = (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[1])) & (InitAccumLoop_1_iacc_6_0_sva_5_0[5]);
  assign and_dcpl_178 = and_dcpl_177 & and_dcpl_176;
  assign and_dcpl_179 = ~((InitAccumLoop_1_iacc_6_0_sva_5_0[3:2]!=2'b00));
  assign and_dcpl_180 = ~((InitAccumLoop_1_iacc_6_0_sva_5_0[0]) | (InitAccumLoop_1_iacc_6_0_sva_5_0[4]));
  assign and_dcpl_181 = and_dcpl_180 & and_dcpl_179;
  assign and_dcpl_185 = IndexLoop_stage_0 & IndexLoop_stage_0_2 & (~ IndexLoop_asn_3_itm_1);
  assign and_dcpl_188 = (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[1:0]==2'b01)
      & IndexLoop_stage_0_2;
  assign and_dcpl_189 = ~((nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[3:2]!=2'b00));
  assign or_dcpl_492 = (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[1:0]!=2'b01);
  assign or_dcpl_493 = (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[3:2]!=2'b00);
  assign or_dcpl_494 = or_dcpl_493 | (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[4]);
  assign or_dcpl_495 = or_dcpl_494 | or_dcpl_492;
  assign and_dcpl_194 = and_dcpl_176 & (~ (ReuseLoop_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_outidx_const_assign_1_ReuseLoop_2_asn_tmp_3_2_0_psp_sva_1[0]));
  assign or_tmp_384 = IndexLoop_asn_3_itm_1 | (~ IndexLoop_stage_0);
  assign mux_487_nl = MUX_s_1_2_2(or_864_cse, (fsm_output[7]), or_888_cse);
  assign mux_tmp_488 = MUX_s_1_2_2((mux_487_nl), or_tmp_48, fsm_output[3]);
  assign and_dcpl_197 = (InitAccumLoop_1_iacc_6_0_sva_5_0[1]) & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[5]))
      & IndexLoop_stage_0_2;
  assign and_dcpl_198 = (InitAccumLoop_1_iacc_6_0_sva_5_0[3:2]==2'b11);
  assign and_dcpl_199 = (InitAccumLoop_1_iacc_6_0_sva_5_0[0]) & (InitAccumLoop_1_iacc_6_0_sva_5_0[4]);
  assign and_dcpl_200 = and_dcpl_199 & and_dcpl_198;
  assign and_dcpl_204 = (~ (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[0]))
      & (~ IndexLoop_stage_0) & IndexLoop_stage_0_2;
  assign and_dcpl_205 = ~((nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[4])
      | (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[1]));
  assign and_dcpl_206 = (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[3:2]==2'b10);
  assign and_dcpl_207 = and_dcpl_206 & and_dcpl_205;
  assign or_dcpl_498 = (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[1:0]!=2'b00);
  assign or_dcpl_499 = (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[3:2]!=2'b10);
  assign or_dcpl_500 = or_dcpl_499 | (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[4]);
  assign or_dcpl_501 = or_dcpl_500 | or_dcpl_498;
  assign and_dcpl_210 = ~(IndexLoop_stage_0 | IndexLoop_stage_0_2);
  assign mux_tmp_496 = MUX_s_1_2_2(or_864_cse, (fsm_output[7]), or_1405_cse);
  assign mux_tmp_497 = MUX_s_1_2_2(mux_509_cse, mux_tmp_496, fsm_output[2]);
  assign mux_tmp_498 = MUX_s_1_2_2(mux_509_cse, mux_tmp_488, fsm_output[2]);
  assign mux_tmp_500 = MUX_s_1_2_2(mux_509_cse, mux_tmp_488, and_817_cse);
  assign and_dcpl_211 = (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[0])) & (InitAccumLoop_1_iacc_6_0_sva_5_0[4]);
  assign and_dcpl_212 = and_dcpl_211 & and_dcpl_198;
  assign and_dcpl_216 = (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[0])
      & (~ IndexLoop_stage_0) & IndexLoop_stage_0_2;
  assign and_dcpl_217 = (~ (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[4]))
      & (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[1]);
  assign and_dcpl_218 = (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[3:2]==2'b01);
  assign and_dcpl_219 = and_dcpl_218 & and_dcpl_217;
  assign or_dcpl_502 = ~((nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[1:0]==2'b11));
  assign or_dcpl_503 = (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[3:2]!=2'b01);
  assign or_dcpl_504 = or_dcpl_503 | (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[4]);
  assign or_dcpl_505 = or_dcpl_504 | or_dcpl_502;
  assign and_dcpl_223 = (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[1])) & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[5]))
      & IndexLoop_stage_0_2;
  assign and_dcpl_227 = (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[1:0]==2'b10)
      & IndexLoop_stage_0_2;
  assign and_dcpl_228 = (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[3:2]==2'b11);
  assign and_dcpl_229 = and_dcpl_228 & (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[4]);
  assign or_dcpl_510 = (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[1:0]!=2'b10);
  assign or_dcpl_511 = ~((nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[3:2]==2'b11));
  assign or_dcpl_512 = or_dcpl_511 | (~ (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[4]));
  assign or_dcpl_513 = or_dcpl_512 | or_dcpl_510;
  assign mux_512_nl = MUX_s_1_2_2(mux_249_cse, or_1213_cse, fsm_output[4]);
  assign mux_tmp_513 = MUX_s_1_2_2((mux_512_nl), or_tmp_48, fsm_output[3]);
  assign mux_tmp_515 = MUX_s_1_2_2(mux_tmp_183, or_1213_cse, fsm_output[4]);
  assign mux_tmp_516 = MUX_s_1_2_2(mux_tmp_515, or_tmp_48, fsm_output[3]);
  assign mux_tmp_517 = MUX_s_1_2_2(mux_tmp_516, mux_tmp_513, fsm_output[2]);
  assign mux_tmp_519 = MUX_s_1_2_2(mux_tmp_184, mux_tmp_513, fsm_output[2]);
  assign mux_tmp_520 = MUX_s_1_2_2(mux_tmp_519, mux_tmp_517, fsm_output[1]);
  assign mux_tmp_521 = MUX_s_1_2_2(mux_tmp_184, mux_tmp_516, fsm_output[2]);
  assign and_dcpl_234 = (InitAccumLoop_1_iacc_6_0_sva_5_0[1]) & (InitAccumLoop_1_iacc_6_0_sva_5_0[5]);
  assign and_dcpl_235 = and_dcpl_234 & IndexLoop_stage_0_2;
  assign and_dcpl_238 = (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[4])
      & (~ (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[1]));
  assign and_dcpl_239 = and_dcpl_218 & and_dcpl_238;
  assign or_dcpl_515 = or_dcpl_503 | (~ (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[4]));
  assign or_dcpl_516 = or_dcpl_515 | or_dcpl_498;
  assign or_dcpl_517 = or_dcpl_512 | or_dcpl_492;
  assign mux_tmp_530 = MUX_s_1_2_2(mux_249_cse, or_1213_cse, or_941_cse);
  assign mux_tmp_532 = MUX_s_1_2_2(or_tmp_196, or_1213_cse, or_941_cse);
  assign and_dcpl_246 = (InitAccumLoop_1_iacc_6_0_sva_5_0[0]) & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[4]));
  assign and_dcpl_247 = and_dcpl_246 & and_dcpl_179;
  assign and_dcpl_250 = (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[4])
      & (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[1]);
  assign and_dcpl_251 = and_dcpl_228 & and_dcpl_250;
  assign and_dcpl_254 = (InitAccumLoop_1_iacc_6_0_sva_5_0[3:2]==2'b10);
  assign and_dcpl_255 = and_dcpl_199 & and_dcpl_254;
  assign or_dcpl_518 = or_dcpl_504 | or_dcpl_510;
  assign mux_540_nl = MUX_s_1_2_2(or_dcpl_334, or_1213_cse, fsm_output[4]);
  assign mux_tmp_541 = MUX_s_1_2_2((mux_540_nl), or_tmp_231, fsm_output[3]);
  assign mux_542_nl = MUX_s_1_2_2(or_tmp_196, or_1213_cse, fsm_output[4]);
  assign mux_tmp_543 = MUX_s_1_2_2((mux_542_nl), or_tmp_231, fsm_output[3]);
  assign and_dcpl_261 = and_dcpl_177 & IndexLoop_stage_0_2;
  assign and_dcpl_262 = (InitAccumLoop_1_iacc_6_0_sva_5_0[3:2]==2'b01);
  assign and_dcpl_263 = and_dcpl_180 & and_dcpl_262;
  assign and_dcpl_266 = and_dcpl_211 & and_dcpl_254;
  assign or_dcpl_519 = or_dcpl_499 | (~ (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[4]));
  assign or_dcpl_520 = or_dcpl_519 | or_dcpl_502;
  assign mux_tmp_549 = MUX_s_1_2_2(or_dcpl_455, or_tmp_231, fsm_output[3]);
  assign mux_tmp_551 = MUX_s_1_2_2(mux_tmp_377, mux_tmp_549, fsm_output[2]);
  assign mux_tmp_552 = MUX_s_1_2_2(or_611_cse, mux_tmp_549, fsm_output[2]);
  assign mux_tmp_553 = MUX_s_1_2_2(mux_tmp_552, mux_tmp_551, fsm_output[1]);
  assign mux_tmp_555 = MUX_s_1_2_2(mux_389_cse, mux_tmp_552, fsm_output[1]);
  assign and_dcpl_274 = and_dcpl_246 & and_dcpl_262;
  assign and_dcpl_277 = and_dcpl_189 & and_dcpl_250;
  assign or_dcpl_521 = or_dcpl_493 | (~ (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[4]));
  assign or_dcpl_522 = or_dcpl_521 | or_dcpl_510;
  assign and_dcpl_283 = and_dcpl_206 & and_dcpl_250;
  assign or_dcpl_525 = or_dcpl_519 | or_dcpl_510;
  assign or_dcpl_526 = or_dcpl_512 | or_dcpl_498;
  assign and_dcpl_295 = and_dcpl_206 & and_dcpl_238;
  assign or_dcpl_528 = or_dcpl_519 | or_dcpl_492;
  assign mux_tmp_570 = MUX_s_1_2_2(mux_tmp_516, mux_509_cse, fsm_output[2]);
  assign or_dcpl_529 = or_dcpl_500 | or_dcpl_492;
  assign and_dcpl_303 = and_dcpl_199 & and_dcpl_262;
  assign or_dcpl_531 = or_dcpl_519 | or_dcpl_498;
  assign and_dcpl_309 = and_dcpl_211 & and_dcpl_262;
  assign and_dcpl_312 = and_dcpl_218 & and_dcpl_250;
  assign or_dcpl_533 = or_dcpl_515 | or_dcpl_502;
  assign or_tmp_449 = (fsm_output[7:3]!=5'b10000);
  assign mux_585_nl = MUX_s_1_2_2(or_611_cse, or_tmp_449, fsm_output[2]);
  assign mux_tmp_586 = MUX_s_1_2_2((mux_585_nl), mux_tmp_552, fsm_output[1]);
  assign mux_tmp_587 = MUX_s_1_2_2(or_611_cse, or_tmp_449, and_817_cse);
  assign or_dcpl_534 = or_dcpl_515 | or_dcpl_510;
  assign mux_tmp_594 = MUX_s_1_2_2(or_611_cse, mux_tmp_549, and_817_cse);
  assign or_dcpl_535 = or_dcpl_515 | or_dcpl_492;
  assign mux_453_nl = MUX_s_1_2_2((fsm_output[2]), (~ (fsm_output[2])), fsm_output[1]);
  assign mux_609_nl = MUX_s_1_2_2(or_10_cse, (mux_453_nl), fsm_output[0]);
  assign and_dcpl_324 = and_dcpl_100 & (mux_609_nl) & (fsm_output[3]);
  assign and_dcpl_325 = and_dcpl_234 & and_dcpl_176;
  assign and_dcpl_326 = and_dcpl_246 & and_dcpl_254;
  assign and_dcpl_329 = and_dcpl_228 & and_dcpl_205;
  assign or_dcpl_536 = or_dcpl_511 | (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[4]);
  assign or_dcpl_537 = or_dcpl_536 | or_dcpl_498;
  assign and_dcpl_334 = and_dcpl_199 & and_dcpl_179;
  assign mux_tmp_620 = MUX_s_1_2_2(mux_tmp_516, mux_tmp_488, fsm_output[2]);
  assign mux_tmp_622 = MUX_s_1_2_2(mux_tmp_570, mux_tmp_620, fsm_output[1]);
  assign and_dcpl_338 = and_dcpl_100 & (and_810_cse_1 ^ (fsm_output[2])) & (fsm_output[3]);
  assign and_dcpl_339 = and_dcpl_180 & and_dcpl_198;
  assign or_dcpl_538 = or_dcpl_536 | or_dcpl_492;
  assign or_dcpl_539 = (ReuseLoop_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_outidx_const_assign_1_ReuseLoop_2_asn_tmp_3_2_0_psp_sva_1[1:0]!=2'b00);
  assign or_dcpl_540 = or_dcpl_539 | (~ (ReuseLoop_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_outidx_const_assign_1_ReuseLoop_2_asn_tmp_3_2_0_psp_sva_1[2]));
  assign and_dcpl_347 = and_dcpl_211 & and_dcpl_179;
  assign or_dcpl_541 = or_dcpl_521 | or_dcpl_502;
  assign mux_tmp_634 = MUX_s_1_2_2(mux_tmp_515, or_tmp_48, or_647_cse_1);
  assign mux_tmp_635 = MUX_s_1_2_2(mux_tmp_620, mux_tmp_634, fsm_output[1]);
  assign and_dcpl_353 = and_dcpl_100 & and_2650_cse & nand_209_cse;
  assign and_dcpl_354 = and_dcpl_246 & and_dcpl_198;
  assign and_dcpl_357 = and_dcpl_228 & and_dcpl_217;
  assign or_dcpl_543 = or_dcpl_536 | or_dcpl_510;
  assign or_dcpl_544 = or_dcpl_539 | (~ nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_out_index_3_0_sva_1_2);
  assign mux_tmp_642 = MUX_s_1_2_2(mux_389_cse, mux_tmp_551, fsm_output[1]);
  assign and_dcpl_365 = and_dcpl_218 & and_dcpl_205;
  assign or_dcpl_545 = or_dcpl_504 | or_dcpl_492;
  assign mux_tmp_646 = MUX_s_1_2_2(mux_tmp_516, mux_tmp_488, and_817_cse);
  assign and_dcpl_369 = and_dcpl_100 & and_2650_cse & ((fsm_output[1]) ^ (fsm_output[0]));
  assign or_dcpl_546 = or_dcpl_536 | or_dcpl_502;
  assign and_dcpl_378 = and_dcpl_189 & and_dcpl_238;
  assign or_dcpl_547 = or_dcpl_521 | or_dcpl_492;
  assign mux_tmp_657 = MUX_s_1_2_2(mux_tmp_517, mux_tmp_634, fsm_output[1]);
  assign or_dcpl_548 = or_dcpl_521 | or_dcpl_498;
  assign mux_tmp_670 = MUX_s_1_2_2(mux_tmp_516, mux_tmp_513, and_817_cse);
  assign mux_tmp_678 = MUX_s_1_2_2(mux_tmp_377, mux_tmp_541, fsm_output[2]);
  assign mux_tmp_679 = MUX_s_1_2_2(mux_tmp_551, mux_tmp_678, fsm_output[1]);
  assign mux_tmp_680 = MUX_s_1_2_2(mux_tmp_377, mux_tmp_549, and_817_cse);
  assign mux_tmp_691 = MUX_s_1_2_2(mux_tmp_377, mux_tmp_541, and_817_cse);
  assign mux_tmp_707 = MUX_s_1_2_2(mux_tmp_521, mux_tmp_517, fsm_output[1]);
  assign and_dcpl_410 = (fsm_output[4:3]==2'b01);
  assign and_dcpl_415 = and_dcpl_189 & and_dcpl_217;
  assign or_dcpl_551 = or_dcpl_494 | or_dcpl_510;
  assign mux_tmp_713 = MUX_s_1_2_2(mux_tmp_377, mux_tmp_543, fsm_output[2]);
  assign mux_tmp_722 = MUX_s_1_2_2(mux_tmp_543, mux_tmp_541, fsm_output[2]);
  assign mux_tmp_723 = MUX_s_1_2_2(mux_tmp_678, mux_tmp_722, fsm_output[1]);
  assign mux_tmp_724 = MUX_s_1_2_2(mux_tmp_713, mux_tmp_678, fsm_output[1]);
  assign and_dcpl_424 = and_dcpl_180 & and_dcpl_254;
  assign and_dcpl_427 = and_dcpl_206 & and_dcpl_217;
  assign or_dcpl_552 = or_dcpl_500 | or_dcpl_502;
  assign and_dcpl_430 = (nand_52_cse | (~ (fsm_output[0]))) & (fsm_output[3]);
  assign mux_tmp_738 = MUX_s_1_2_2(mux_tmp_713, mux_tmp_722, fsm_output[1]);
  assign or_dcpl_554 = or_dcpl_500 | or_dcpl_510;
  assign mux_tmp_742 = MUX_s_1_2_2(mux_tmp_184, mux_tmp_530, fsm_output[2]);
  assign and_dcpl_449 = nor_298_cse & and_dcpl_73 & (fsm_output[0]) & (~ IndexLoop_stage_0)
      & IndexLoop_stage_0_2;
  assign mux_tmp_771 = MUX_s_1_2_2(or_dcpl_334, or_1213_cse, or_941_cse);
  assign mux_tmp_772 = MUX_s_1_2_2(mux_tmp_543, mux_tmp_771, fsm_output[2]);
  assign mux_tmp_773 = MUX_s_1_2_2(mux_tmp_722, mux_tmp_772, fsm_output[1]);
  assign mux_tmp_774 = MUX_s_1_2_2(mux_tmp_543, mux_tmp_541, and_817_cse);
  assign or_dcpl_556 = or_dcpl_504 | or_dcpl_498;
  assign and_dcpl_467 = and_dcpl_100 & and_dcpl_430;
  assign mux_tmp_787 = MUX_s_1_2_2(mux_tmp_543, mux_tmp_771, and_817_cse);
  assign mux_tmp_806 = MUX_s_1_2_2(mux_tmp_532, mux_tmp_184, fsm_output[2]);
  assign mux_tmp_814 = MUX_s_1_2_2(mux_tmp_543, mux_tmp_532, fsm_output[2]);
  assign mux_tmp_819 = MUX_s_1_2_2(mux_tmp_532, mux_tmp_530, fsm_output[2]);
  assign mux_tmp_820 = MUX_s_1_2_2(mux_tmp_819, mux_tmp_742, fsm_output[1]);
  assign and_dcpl_486 = and_dcpl_228 & and_dcpl_238;
  assign mux_tmp_829 = MUX_s_1_2_2(mux_tmp_532, mux_tmp_771, fsm_output[2]);
  assign mux_tmp_830 = MUX_s_1_2_2(mux_tmp_772, mux_tmp_829, fsm_output[1]);
  assign mux_tmp_831 = MUX_s_1_2_2(mux_tmp_814, mux_tmp_772, fsm_output[1]);
  assign mux_tmp_837 = MUX_s_1_2_2(mux_tmp_806, mux_tmp_819, fsm_output[1]);
  assign mux_tmp_845 = MUX_s_1_2_2(mux_tmp_814, mux_tmp_829, fsm_output[1]);
  assign or_dcpl_558 = or_dcpl_494 | or_dcpl_502;
  assign mux_tmp_860 = MUX_s_1_2_2(mux_tmp_829, mux_tmp_819, fsm_output[1]);
  assign mux_tmp_861 = MUX_s_1_2_2(mux_tmp_532, mux_tmp_530, and_817_cse);
  assign or_dcpl_559 = or_dcpl_512 | or_dcpl_502;
  assign mux_tmp_870 = MUX_s_1_2_2(mux_tmp_532, mux_tmp_771, and_817_cse);
  assign and_dcpl_509 = and_dcpl_189 & and_dcpl_205;
  assign or_dcpl_560 = or_dcpl_376 | or_dcpl_363;
  assign or_dcpl_561 = or_dcpl_494 | or_dcpl_498;
  assign and_dcpl_517 = and_2650_cse & and_dcpl_103;
  assign and_dcpl_519 = and_dcpl_171 & nor_306_cse;
  assign and_dcpl_520 = and_dcpl_54 & and_dcpl_519;
  assign or_1391_nl = (fsm_output[6:3]!=4'b0000);
  assign mux_tmp_909 = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), or_1391_nl);
  assign mux_tmp_911 = MUX_s_1_2_2(mux_tmp_909, mux_tmp_496, and_817_cse);
  assign or_dcpl_571 = or_dcpl_376 | or_dcpl_362;
  assign or_dcpl_572 = or_dcpl_381 | or_dcpl_368;
  assign or_dcpl_573 = or_dcpl_365 | or_dcpl_362;
  assign or_dcpl_574 = or_dcpl_371 | or_dcpl_368;
  assign or_dcpl_575 = or_dcpl_376 | or_dcpl_373;
  assign or_dcpl_576 = or_dcpl_381 | or_dcpl_378;
  assign or_dcpl_577 = or_dcpl_365 | or_dcpl_373;
  assign or_dcpl_578 = or_dcpl_371 | or_dcpl_378;
  assign or_dcpl_579 = or_dcpl_376 | or_dcpl_378;
  assign or_dcpl_580 = or_dcpl_381 | or_dcpl_373;
  assign or_dcpl_581 = or_dcpl_365 | or_dcpl_378;
  assign or_dcpl_582 = or_dcpl_371 | or_dcpl_373;
  assign or_dcpl_583 = or_dcpl_376 | or_dcpl_368;
  assign or_dcpl_584 = or_dcpl_381 | or_dcpl_362;
  assign or_dcpl_585 = or_dcpl_365 | or_dcpl_368;
  assign or_dcpl_586 = or_dcpl_371 | or_dcpl_362;
  assign or_dcpl_587 = or_dcpl_397 | or_dcpl_362;
  assign or_dcpl_588 = or_dcpl_399 | or_dcpl_368;
  assign or_dcpl_589 = or_dcpl_401 | or_dcpl_362;
  assign or_dcpl_590 = or_dcpl_403 | or_dcpl_368;
  assign or_dcpl_591 = or_dcpl_397 | or_dcpl_373;
  assign or_dcpl_592 = or_dcpl_399 | or_dcpl_378;
  assign or_dcpl_593 = or_dcpl_401 | or_dcpl_373;
  assign or_dcpl_594 = or_dcpl_403 | or_dcpl_378;
  assign or_dcpl_595 = or_dcpl_397 | or_dcpl_378;
  assign or_dcpl_596 = or_dcpl_399 | or_dcpl_373;
  assign or_dcpl_597 = or_dcpl_401 | or_dcpl_378;
  assign or_dcpl_598 = or_dcpl_403 | or_dcpl_373;
  assign or_dcpl_599 = or_dcpl_397 | or_dcpl_368;
  assign or_dcpl_600 = or_dcpl_399 | or_dcpl_362;
  assign or_dcpl_601 = or_dcpl_401 | or_dcpl_368;
  assign or_dcpl_602 = or_dcpl_403 | or_dcpl_362;
  assign mux_tmp_913 = MUX_s_1_2_2((fsm_output[6]), or_tmp_91, or_1405_cse);
  assign mux_tmp_914 = MUX_s_1_2_2(or_865_cse_1, or_tmp_91, or_1405_cse);
  assign mux_tmp_915 = MUX_s_1_2_2(mux_tmp_914, mux_tmp_913, fsm_output[2]);
  assign mux_tmp_918 = MUX_s_1_2_2(mux_tmp_914, mux_tmp_913, and_817_cse);
  assign mux_tmp_925 = MUX_s_1_2_2(mux_509_cse, mux_tmp_909, fsm_output[2]);
  assign mux_924_nl = MUX_s_1_2_2(mux_tmp_909, mux_tmp_496, fsm_output[2]);
  assign mux_tmp_926 = MUX_s_1_2_2(mux_tmp_925, (mux_924_nl), fsm_output[1]);
  assign and_dcpl_567 = and_dcpl_171 & and_dcpl_56;
  assign and_dcpl_570 = and_dcpl_171 & and_dcpl_103;
  assign mux_tmp_928 = MUX_s_1_2_2(mux_tmp_925, mux_tmp_497, fsm_output[1]);
  assign and_dcpl_573 = and_dcpl_171 & and_810_cse_1;
  assign and_dcpl_576 = and_2650_cse & nor_306_cse;
  assign mux_tmp_930 = MUX_s_1_2_2(mux_509_cse, mux_tmp_496, and_817_cse);
  assign and_dcpl_579 = and_2650_cse & and_dcpl_56;
  assign and_dcpl_584 = and_2650_cse & and_810_cse_1;
  assign and_dcpl_587 = nor_942_cse & nor_306_cse;
  assign and_dcpl_588 = nor_944_cse & and_dcpl_99;
  assign mux_tmp_933 = MUX_s_1_2_2(mux_tmp_570, mux_tmp_498, fsm_output[1]);
  assign and_dcpl_590 = and_dcpl_58 & and_dcpl_99;
  assign and_dcpl_592 = nor_942_cse & and_dcpl_56;
  assign and_dcpl_623 = (fsm_output[5:4]==2'b10);
  assign and_dcpl_624 = nor_944_cse & and_dcpl_623;
  assign and_dcpl_626 = and_dcpl_58 & and_dcpl_623;
  assign and_dcpl_658 = (fsm_output[5:4]==2'b11);
  assign and_dcpl_659 = nor_944_cse & and_dcpl_658;
  assign and_dcpl_661 = and_dcpl_58 & and_dcpl_658;
  assign or_dcpl_607 = (fsm_output[3:2]!=2'b10);
  assign or_dcpl_611 = (fsm_output[1:0]!=2'b01);
  assign layer7_out_rsci_idat_11_0_mx0c1 = and_dcpl_87 & and_dcpl_84 & IndexLoop_stage_0
      & (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_1_or_tmp);
  assign layer7_out_rsci_idat_29_18_mx0c1 = or_dcpl_339 & and_dcpl_70 & and_dcpl_106;
  assign layer7_out_rsci_idat_47_36_mx0c1 = or_dcpl_341 & and_dcpl_70 & and_dcpl_106;
  assign layer7_out_rsci_idat_65_54_mx0c1 = or_dcpl_343 & and_dcpl_70 & and_dcpl_106;
  assign layer7_out_rsci_idat_83_72_mx0c1 = or_dcpl_346 & and_dcpl_70 & and_dcpl_106;
  assign layer7_out_rsci_idat_101_90_mx0c1 = or_dcpl_347 & and_dcpl_70 & and_dcpl_106;
  assign layer7_out_rsci_idat_119_108_mx0c1 = or_dcpl_348 & and_dcpl_70 & and_dcpl_106;
  assign layer7_out_rsci_idat_137_126_mx0c1 = or_dcpl_349 & and_dcpl_70 & and_dcpl_106;
  assign layer7_out_rsci_idat_155_144_mx0c1 = or_dcpl_351 & and_dcpl_70 & and_dcpl_106;
  assign layer7_out_rsci_idat_173_162_mx0c1 = (or_dcpl_350 | or_dcpl_337) & and_dcpl_70
      & and_dcpl_106;
  assign mux_491_itm = MUX_s_1_2_2(mux_509_cse, mux_tmp_488, and_2657_cse);
  assign mux_499_nl = MUX_s_1_2_2(mux_tmp_498, mux_tmp_497, fsm_output[1]);
  assign mux_501_itm = MUX_s_1_2_2(mux_tmp_500, (mux_499_nl), fsm_output[0]);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_sva_2_mx0c3
      = and_dcpl_54 & (nor_306_cse | (~ (fsm_output[2]))) & (fsm_output[3]);
  assign mux_533_itm = MUX_s_1_2_2(mux_tmp_532, mux_tmp_530, and_2657_cse);
  assign mux_544_itm = MUX_s_1_2_2(mux_tmp_543, mux_tmp_541, and_2657_cse);
  assign mux_556_itm = MUX_s_1_2_2(mux_tmp_555, mux_tmp_553, fsm_output[0]);
  assign mux_563_nl = MUX_s_1_2_2(mux_425_cse, mux_421_cse, fsm_output[0]);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_sva_2_mx0c2
      = (~ (mux_563_nl)) & and_dcpl_169;
  assign mux_568_nl = MUX_s_1_2_2(mux_tmp_419, mux_421_cse, fsm_output[0]);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_sva_2_mx0c2
      = (~ (mux_568_nl)) & and_dcpl_169;
  assign mux_571_itm = MUX_s_1_2_2(mux_tmp_570, mux_tmp_498, or_1875_cse);
  assign mux_579_nl = MUX_s_1_2_2(nand_tmp_14, mux_33_cse, or_1875_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_sva_2_mx0c2
      = (~ (mux_579_nl)) & and_dcpl_169;
  assign mux_582_nl = MUX_s_1_2_2(mux_661_cse, or_864_cse, and_2657_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_sva_2_mx0c2
      = (~ (mux_582_nl)) & and_dcpl_169;
  assign mux_588_itm = MUX_s_1_2_2(mux_tmp_587, mux_tmp_586, fsm_output[0]);
  assign mux_595_itm = MUX_s_1_2_2(mux_tmp_594, mux_tmp_586, fsm_output[0]);
  assign mux_616_itm = MUX_s_1_2_2(or_611_cse, mux_tmp_549, and_2657_cse);
  assign mux_631_itm = MUX_s_1_2_2(mux_389_cse, mux_tmp_552, or_1875_cse);
  assign mux_643_itm = MUX_s_1_2_2(mux_tmp_642, mux_tmp_553, fsm_output[0]);
  assign mux_654_itm = MUX_s_1_2_2(mux_389_cse, mux_tmp_551, or_1875_cse);
  assign mux_665_itm = MUX_s_1_2_2(mux_tmp_377, mux_tmp_549, and_2657_cse);
  assign mux_681_itm = MUX_s_1_2_2(mux_tmp_680, mux_tmp_679, fsm_output[0]);
  assign mux_692_itm = MUX_s_1_2_2(mux_tmp_691, mux_tmp_679, fsm_output[0]);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_sva_2_mx0c3
      = and_dcpl_54 & and_dcpl_171 & nand_209_cse;
  assign mux_703_itm = MUX_s_1_2_2(mux_tmp_377, mux_tmp_541, and_2657_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_sva_2_mx0c3
      = and_dcpl_70 & and_dcpl_410 & (~ (fsm_output[2]));
  assign mux_714_itm = MUX_s_1_2_2(mux_tmp_713, mux_tmp_678, or_1875_cse);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_sva_2_mx0c3
      = and_dcpl_54 & nand_52_cse & (fsm_output[3]);
  assign mux_725_itm = MUX_s_1_2_2(mux_tmp_724, mux_tmp_723, fsm_output[0]);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_sva_2_mx0c3
      = and_dcpl_54 & and_dcpl_430;
  assign mux_739_itm = MUX_s_1_2_2(mux_tmp_738, mux_tmp_723, fsm_output[0]);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_sva_2_mx0c3
      = and_dcpl_70 & and_dcpl_410;
  assign mux_753_itm = MUX_s_1_2_2(mux_tmp_713, mux_tmp_722, or_1875_cse);
  assign mux_3_nl = MUX_s_1_2_2(mux_tmp_2, or_tmp_1, fsm_output[2]);
  assign mux_1_nl = MUX_s_1_2_2(mux_cse, or_tmp_1, fsm_output[2]);
  assign mux_4_nl = MUX_s_1_2_2((mux_3_nl), (mux_1_nl), fsm_output[1]);
  assign mux_761_nl = MUX_s_1_2_2((mux_4_nl), or_tmp_1, fsm_output[0]);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_2_mx0c0
      = (~ (mux_761_nl)) & and_dcpl;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_2_mx0c3
      = or_dcpl_531 & and_dcpl_75 & and_dcpl_449;
  assign or_867_nl = (~ (fsm_output[1])) | (fsm_output[6]) | (~ (fsm_output[7]));
  assign mux_481_nl = MUX_s_1_2_2(or_865_cse_1, or_864_cse, fsm_output[1]);
  assign mux_762_nl = MUX_s_1_2_2((or_867_nl), (mux_481_nl), IndexLoop_stage_0);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_2_mx0c4
      = (~ (mux_762_nl)) & (~ (fsm_output[5])) & nor_298_cse & (fsm_output[2]) &
      (fsm_output[0]);
  assign mux_764_nl = MUX_s_1_2_2(nor_942_cse, mux_456_cse, and_810_cse_1);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_2_mx0c5
      = (~ (mux_764_nl)) & and_dcpl_100;
  assign mux_775_itm = MUX_s_1_2_2(mux_tmp_774, mux_tmp_773, fsm_output[0]);
  assign or_11_nl = (fsm_output[3]) | (fsm_output[7]);
  assign mux_8_nl = MUX_s_1_2_2(nand_198_cse, (or_11_nl), fsm_output[1]);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_2_mx0c0
      = ~((mux_8_nl) | (fsm_output[6]) | (~ nor_943_cse) | (fsm_output[2]) | (fsm_output[0]));
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_2_mx0c4
      = and_dcpl_54 & and_dcpl_50 & (fsm_output[1]);
  assign mux_788_itm = MUX_s_1_2_2(mux_tmp_787, mux_tmp_773, fsm_output[0]);
  assign mux_802_itm = MUX_s_1_2_2(mux_tmp_543, mux_tmp_771, and_2657_cse);
  assign mux_815_itm = MUX_s_1_2_2(mux_tmp_814, mux_tmp_772, or_1875_cse);
  assign mux_832_itm = MUX_s_1_2_2(mux_tmp_831, mux_tmp_830, fsm_output[0]);
  assign mux_846_itm = MUX_s_1_2_2(mux_tmp_845, mux_tmp_830, fsm_output[0]);
  assign mux_850_itm = MUX_s_1_2_2(mux_tmp_806, mux_tmp_819, or_1875_cse);
  assign mux_856_itm = MUX_s_1_2_2(mux_tmp_814, mux_tmp_829, or_1875_cse);
  assign mux_862_itm = MUX_s_1_2_2(mux_tmp_861, mux_tmp_860, fsm_output[0]);
  assign mux_867_itm = MUX_s_1_2_2(mux_tmp_532, mux_tmp_771, and_2657_cse);
  assign mux_872_itm = MUX_s_1_2_2(mux_tmp_870, mux_tmp_860, fsm_output[0]);
  assign MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_mx0c2
      = or_dcpl_427 & nor_944_cse & nor_943_cse & nor_942_cse & and_810_cse_1 & and_dcpl_176;
  assign MultLoop_2_and_28_m1c = (ROM_1i9_1o3_2fa806bf16b3e0d54016201674d036b62f_1==3'b001)
      & IndexLoop_stage_0;
  assign MultLoop_2_and_29_m1c = (ROM_1i9_1o3_2fa806bf16b3e0d54016201674d036b62f_1==3'b010)
      & IndexLoop_stage_0;
  assign MultLoop_2_and_30_m1c = (ROM_1i9_1o3_2fa806bf16b3e0d54016201674d036b62f_1==3'b011)
      & IndexLoop_stage_0;
  assign MultLoop_2_and_31_m1c = (ROM_1i9_1o3_2fa806bf16b3e0d54016201674d036b62f_1==3'b100)
      & IndexLoop_stage_0;
  assign MultLoop_2_and_26_m1c = (~ or_1479_cse) & MultLoop_2_nor_m1c & IndexLoop_stage_0;
  assign MultLoop_2_and_m1c = (MultLoop_2_1_acc_3_tmp==3'b001);
  assign and_550_m1c = or_dcpl_445 & and_dcpl_176;
  assign MultLoop_2_and_21_m1c = (~ or_1479_cse) & MultLoop_2_and_m1c & IndexLoop_stage_0;
  assign MultLoop_2_and_20_m1c = (MultLoop_2_1_acc_3_tmp==3'b000) & IndexLoop_stage_0;
  assign MultLoop_2_and_25_m1c = (MultLoop_2_1_acc_3_tmp==3'b111) & IndexLoop_stage_0;
  assign MultLoop_2_and_24_m1c = (MultLoop_2_1_acc_3_tmp==3'b110) & IndexLoop_stage_0;
  assign MultLoop_2_and_23_m1c = (MultLoop_2_1_acc_3_tmp==3'b101) & IndexLoop_stage_0;
  assign w2_rsci_adra_d = w2_rsci_adra_d_reg;
  assign w2_rsci_ena_d = w2_rsci_ena_d_reg;
  assign w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign w4_rsci_adra_d = w4_rsci_adra_d_reg;
  assign w4_rsci_ena_d = w4_rsci_ena_d_reg;
  assign w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign w6_rsci_adra_d = w6_rsci_adra_d_reg;
  assign w6_rsci_ena_d = w6_rsci_ena_d_reg;
  assign w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign nor_450_nl = ~((fsm_output[7:6]!=2'b01));
  assign mux_988_nl = MUX_s_1_2_2((nor_450_nl), nor_586_cse, fsm_output[1]);
  assign and_dcpl_730 = (mux_988_nl) & (~ (fsm_output[5])) & (~ (fsm_output[4]))
      & (~ (fsm_output[3])) & (fsm_output[2]) & (fsm_output[0]);
  assign and_dcpl_737 = (fsm_output[7:6]==2'b00) & nor_943_cse & (fsm_output[3:0]==4'b0011);
  assign nand_152_cse = ~((fsm_output[2]) & (fsm_output[6]));
  assign mux_966_nl = MUX_s_1_2_2(nand_152_cse, or_1800_cse, fsm_output[1]);
  assign and_dcpl_741 = ~((mux_966_nl) | (fsm_output[7]) | (~ nor_943_cse) | (fsm_output[3])
      | (fsm_output[0]));
  assign and_dcpl_756 = (fsm_output[3:2]==2'b00) & and_810_cse_1;
  assign and_dcpl_760 = and_dcpl_53 & (fsm_output[5:4]==2'b01) & and_dcpl_756;
  assign and_dcpl_764 = (fsm_output[7:6]==2'b00) & nor_943_cse & and_dcpl_756;
  assign and_dcpl_768 = and_dcpl_53 & nor_943_cse & (fsm_output[3:2]==2'b01) & and_810_cse_1;
  assign and_dcpl_779 = (fsm_output[7:4]==4'b0000) & nor_942_cse & (fsm_output[1:0]==2'b11);
  assign and_dcpl_926 = and_dcpl_53 & (fsm_output[5:4]==2'b00);
  assign and_dcpl_949 = and_dcpl_53 & (fsm_output[5:4]==2'b01);
  assign and_1134_cse = and_dcpl_949 & nor_942_cse & and_dcpl_103;
  assign and_dcpl_964 = and_dcpl_53 & (fsm_output[5:2]==4'b0011) & and_dcpl_103;
  assign and_dcpl_967 = and_dcpl_949 & nor_942_cse & (fsm_output[1:0]==2'b11);
  assign and_dcpl_979 = (fsm_output[7:6]==2'b10) & nor_943_cse & (fsm_output[3:0]==4'b0111);
  assign and_1161_cse = (fsm_output[7:6]==2'b00) & nor_943_cse & nor_942_cse & and_810_cse_1;
  assign and_dcpl_992 = (fsm_output[7:6]==2'b01) & nor_943_cse & (fsm_output[3:2]==2'b01)
      & and_dcpl_56;
  assign and_1173_cse = and_dcpl_54 & and_dcpl_171 & nor_306_cse;
  assign and_1175_cse = and_dcpl_54 & and_dcpl_171 & and_dcpl_56;
  assign and_1178_cse = and_dcpl_54 & and_dcpl_171 & and_dcpl_103;
  assign and_1180_cse = and_dcpl_54 & and_dcpl_171 & and_810_cse_1;
  assign and_1183_cse = and_dcpl_54 & and_2650_cse & nor_306_cse;
  assign and_1185_cse = and_dcpl_54 & and_2650_cse & and_dcpl_56;
  assign and_1187_cse = and_dcpl_54 & and_2650_cse & and_dcpl_103;
  assign and_1189_cse = and_dcpl_54 & and_2650_cse & and_810_cse_1;
  assign and_1193_cse = and_dcpl_949 & nor_942_cse & nor_306_cse;
  assign and_1195_cse = and_dcpl_949 & nor_942_cse & and_dcpl_56;
  assign and_1270_cse = and_dcpl_926 & and_dcpl_171 & nor_306_cse;
  assign and_1273_cse = and_dcpl_926 & and_dcpl_171 & and_dcpl_56;
  assign and_1276_cse = and_dcpl_926 & and_dcpl_171 & and_dcpl_103;
  assign and_1279_cse = and_dcpl_926 & and_dcpl_171 & and_810_cse_1;
  assign and_1282_cse = and_dcpl_926 & and_2650_cse & nor_306_cse;
  assign and_1284_cse = and_dcpl_926 & and_2650_cse & and_dcpl_56;
  assign and_1286_cse = and_dcpl_926 & and_2650_cse & and_dcpl_103;
  assign and_1288_cse = and_dcpl_926 & and_2650_cse & and_810_cse_1;
  assign and_dcpl_1163 = (fsm_output[7:4]==4'b1001) & nor_942_cse & (fsm_output[1:0]==2'b11);
  assign and_dcpl_1170 = (fsm_output[7:6]==2'b01) & nor_943_cse & and_dcpl_57;
  assign and_dcpl_1175 = and_dcpl_53 & nor_943_cse & and_dcpl_51;
  assign and_dcpl_1180 = and_dcpl_949 & and_dcpl_50 & nor_306_cse;
  assign and_dcpl_1181 = and_dcpl_949 & and_dcpl_57;
  assign and_dcpl_1184 = and_dcpl_949 & and_dcpl_50 & and_dcpl_103;
  assign and_dcpl_1185 = and_dcpl_949 & and_dcpl_51;
  assign and_dcpl_1188 = and_dcpl_949 & and_dcpl_171 & nor_306_cse;
  assign and_dcpl_1190 = and_dcpl_949 & and_dcpl_171 & and_dcpl_56;
  assign and_dcpl_1192 = and_dcpl_949 & and_dcpl_171 & and_dcpl_103;
  assign and_dcpl_1194 = and_dcpl_949 & and_dcpl_171 & and_810_cse_1;
  assign and_dcpl_1197 = and_dcpl_949 & and_2650_cse & nor_306_cse;
  assign and_dcpl_1199 = and_dcpl_949 & and_2650_cse & and_dcpl_56;
  assign and_dcpl_1224 = (fsm_output[7:6]==2'b01) & nor_943_cse & and_dcpl_50 & (fsm_output[1:0]==2'b01);
  assign and_dcpl_1228 = (fsm_output[7:6]==2'b10) & nor_943_cse & and_dcpl_50 & and_810_cse_1;
  assign and_dcpl_1278 = ~(((fsm_output[6]) ^ (fsm_output[0])) | (fsm_output[7]));
  assign and_dcpl_1283 = and_dcpl_169 & and_817_cse & and_dcpl_1278;
  assign and_dcpl_1285 = (~ (fsm_output[4])) & (fsm_output[2]);
  assign and_dcpl_1287 = ~((fsm_output[7]) | (fsm_output[5]));
  assign and_dcpl_1289 = and_dcpl_1287 & ((fsm_output[6]) ^ (fsm_output[3])) & and_dcpl_1285
      & and_dcpl_103;
  assign nor_tmp_215 = (fsm_output[3]) & (fsm_output[6]);
  assign nor_441_nl = ~((fsm_output[3]) | (fsm_output[6]));
  assign mux_967_nl = MUX_s_1_2_2((nor_441_nl), nor_tmp_215, fsm_output[1]);
  assign and_dcpl_1293 = (mux_967_nl) & (~ (fsm_output[7])) & nor_943_cse & (fsm_output[2])
      & (~ (fsm_output[0]));
  assign and_dcpl_1294 = (fsm_output[2]) & (fsm_output[0]);
  assign nor_439_nl = ~((fsm_output[3]) | (~ (fsm_output[7])));
  assign nor_440_nl = ~((~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_968_nl = MUX_s_1_2_2((nor_439_nl), (nor_440_nl), fsm_output[1]);
  assign and_dcpl_1297 = (mux_968_nl) & (~ (fsm_output[6])) & nor_943_cse & and_dcpl_1294;
  assign and_dcpl_1301 = and_dcpl_1287 & (~((fsm_output[6]) ^ (fsm_output[3]))) &
      and_dcpl_1285 & and_dcpl_56;
  assign nor_437_nl = ~((fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[6]) |
      (~ (fsm_output[7])));
  assign nor_438_nl = ~((~ (fsm_output[1])) | (fsm_output[2]) | (~ (fsm_output[6]))
      | (fsm_output[7]));
  assign mux_969_nl = MUX_s_1_2_2((nor_437_nl), (nor_438_nl), fsm_output[0]);
  assign and_dcpl_1302 = (mux_969_nl) & and_dcpl_169;
  assign nor_tmp_216 = (fsm_output[4]) & (fsm_output[6]);
  assign nor_435_nl = ~((fsm_output[2:1]!=2'b00) | (~ nor_tmp_216));
  assign nor_436_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[2])) | (fsm_output[4])
      | (fsm_output[6]));
  assign mux_970_nl = MUX_s_1_2_2((nor_435_nl), (nor_436_nl), fsm_output[0]);
  assign and_dcpl_1304 = (mux_970_nl) & and_dcpl_1287 & (~ (fsm_output[3]));
  assign and_dcpl_1306 = (~ (fsm_output[5])) & (fsm_output[3]);
  assign nor_434_nl = ~((fsm_output[4]) | (fsm_output[6]));
  assign mux_971_nl = MUX_s_1_2_2((nor_434_nl), nor_tmp_216, fsm_output[1]);
  assign and_dcpl_1309 = (mux_971_nl) & (~ (fsm_output[7])) & and_dcpl_1306 & (~
      (fsm_output[2])) & (~ (fsm_output[0]));
  assign nor_432_nl = ~((fsm_output[4]) | (~ (fsm_output[6])));
  assign nor_433_nl = ~((~ (fsm_output[4])) | (fsm_output[6]));
  assign mux_972_nl = MUX_s_1_2_2((nor_432_nl), (nor_433_nl), fsm_output[0]);
  assign and_dcpl_1313 = (mux_972_nl) & (~ (fsm_output[7])) & and_dcpl_1306 & nor_668_cse;
  assign and_dcpl_1314 = ~((fsm_output[7]) | (fsm_output[4]));
  assign nor_tmp_217 = (fsm_output[6:5]==2'b11);
  assign nor_430_nl = ~((fsm_output[3:2]!=2'b01) | (~ nor_tmp_217));
  assign nor_431_nl = ~((fsm_output[2]) | (~ (fsm_output[3])) | (fsm_output[5]) |
      (fsm_output[6]));
  assign mux_973_nl = MUX_s_1_2_2((nor_430_nl), (nor_431_nl), fsm_output[0]);
  assign and_dcpl_1316 = (mux_973_nl) & and_dcpl_1314 & (~ (fsm_output[1]));
  assign nor_428_nl = ~((~ (fsm_output[3])) | (fsm_output[5]) | (~ (fsm_output[6])));
  assign nor_429_nl = ~((fsm_output[3]) | (~ (fsm_output[5])) | (fsm_output[6]));
  assign mux_974_nl = MUX_s_1_2_2((nor_428_nl), (nor_429_nl), fsm_output[1]);
  assign and_dcpl_1319 = (mux_974_nl) & and_dcpl_1314 & (~ (fsm_output[2])) & (fsm_output[0]);
  assign mux_975_nl = MUX_s_1_2_2(and_dcpl, nor_tmp_217, fsm_output[2]);
  assign and_dcpl_1323 = (mux_975_nl) & (~ (fsm_output[7])) & and_dcpl_410 & and_dcpl_103;
  assign nor_425_nl = ~((~ (fsm_output[1])) | (fsm_output[2]) | (fsm_output[5]) |
      (~ (fsm_output[6])));
  assign nor_426_nl = ~((fsm_output[1]) | (~ (fsm_output[2])) | (~ (fsm_output[5]))
      | (fsm_output[6]));
  assign mux_976_nl = MUX_s_1_2_2((nor_425_nl), (nor_426_nl), fsm_output[0]);
  assign and_dcpl_1325 = (mux_976_nl) & and_dcpl_1314 & (fsm_output[3]);
  assign nor_423_nl = ~((fsm_output[1]) | (~((fsm_output[6:4]==3'b111))));
  assign nor_424_nl = ~((~ (fsm_output[1])) | (fsm_output[4]) | (fsm_output[5]) |
      (fsm_output[6]));
  assign mux_977_nl = MUX_s_1_2_2((nor_423_nl), (nor_424_nl), fsm_output[0]);
  assign and_dcpl_1328 = (mux_977_nl) & (~ (fsm_output[7])) & (fsm_output[3]) & (~
      (fsm_output[2]));
  assign nor_421_nl = ~((fsm_output[6:3]!=4'b1001));
  assign nor_422_nl = ~((fsm_output[6:3]!=4'b0110));
  assign mux_978_nl = MUX_s_1_2_2((nor_421_nl), (nor_422_nl), fsm_output[2]);
  assign and_dcpl_1331 = (mux_978_nl) & (~ (fsm_output[7])) & (fsm_output[1]) & (fsm_output[0]);
  assign nor_419_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[7]));
  assign nor_420_nl = ~((fsm_output[2]) | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_979_nl = MUX_s_1_2_2((nor_419_nl), (nor_420_nl), fsm_output[1]);
  assign and_dcpl_1334 = (mux_979_nl) & and_dcpl & (~ (fsm_output[4])) & (~ (fsm_output[0]));
  assign mux_980_nl = MUX_s_1_2_2(and_2650_cse, nor_942_cse, fsm_output[0]);
  assign and_dcpl_1339 = (mux_980_nl) & (~ (fsm_output[7])) & (fsm_output[6]) & (~
      (fsm_output[5])) & (~ (fsm_output[4])) & (~ (fsm_output[1]));
  assign and_dcpl_1342 = and_dcpl_1287 & (~((fsm_output[6]) ^ (fsm_output[1]))) &
      and_dcpl_410 & and_dcpl_1294;
  assign and_dcpl_1344 = and_dcpl_99 & (~ (fsm_output[3]));
  assign and_dcpl_1346 = and_dcpl_1344 & nor_668_cse & and_dcpl_1278;
  assign nand_150_nl = ~((fsm_output[1]) & (fsm_output[6]));
  assign or_1473_nl = (fsm_output[1]) | (fsm_output[6]);
  assign mux_981_nl = MUX_s_1_2_2((nand_150_nl), (or_1473_nl), fsm_output[0]);
  assign and_dcpl_1349 = ~((mux_981_nl) | (fsm_output[7]));
  assign and_dcpl_1350 = and_dcpl_1349 & and_dcpl_99 & nor_942_cse;
  assign and_dcpl_1351 = (fsm_output[2:1]==2'b01);
  assign and_dcpl_1353 = and_dcpl_1344 & and_dcpl_1351 & and_dcpl_1278;
  assign and_dcpl_1354 = (fsm_output[4:3]==2'b10);
  assign nor_415_nl = ~((fsm_output[1]) | nand_152_cse);
  assign nor_416_nl = ~((~ (fsm_output[1])) | (fsm_output[2]) | (fsm_output[6]));
  assign not_tmp_680 = MUX_s_1_2_2((nor_415_nl), (nor_416_nl), fsm_output[0]);
  assign and_dcpl_1356 = not_tmp_680 & and_dcpl_1287 & and_dcpl_1354;
  assign and_dcpl_1359 = and_dcpl_1344 & and_dcpl_73 & and_dcpl_1278;
  assign and_dcpl_1362 = and_dcpl_1349 & and_dcpl_99 & and_dcpl_50;
  assign and_dcpl_1364 = and_dcpl_1344 & and_817_cse & and_dcpl_1278;
  assign nor_413_nl = ~((fsm_output[2:1]!=2'b00) | (~ nor_tmp_215));
  assign nor_414_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[2])) | (fsm_output[3])
      | (fsm_output[6]));
  assign not_tmp_682 = MUX_s_1_2_2((nor_413_nl), (nor_414_nl), fsm_output[0]);
  assign and_dcpl_1366 = not_tmp_682 & and_dcpl_1287 & (fsm_output[4]);
  assign and_dcpl_1367 = and_dcpl_99 & (fsm_output[3]);
  assign and_dcpl_1369 = and_dcpl_1367 & nor_668_cse & and_dcpl_1278;
  assign and_dcpl_1371 = and_dcpl_1367 & and_dcpl_1351 & and_dcpl_1278;
  assign and_dcpl_1374 = not_tmp_680 & and_dcpl_1287 & and_862_cse;
  assign and_dcpl_1376 = and_dcpl_1367 & and_dcpl_73 & and_dcpl_1278;
  assign and_dcpl_1378 = and_dcpl_1349 & and_dcpl_99 & and_2650_cse;
  assign and_dcpl_1380 = and_dcpl_1367 & and_817_cse & and_dcpl_1278;
  assign or_nl = (fsm_output[4:1]!=4'b0000) | (~ nor_tmp_217);
  assign or_1472_nl = (fsm_output[6:1]!=6'b001111);
  assign mux_984_nl = MUX_s_1_2_2((or_nl), (or_1472_nl), fsm_output[0]);
  assign and_dcpl_1381 = ~((mux_984_nl) | (fsm_output[7]));
  assign and_dcpl_1383 = and_dcpl_623 & (~ (fsm_output[3]));
  assign and_dcpl_1385 = and_dcpl_1383 & nor_668_cse & and_dcpl_1278;
  assign and_dcpl_1387 = and_dcpl_1349 & and_dcpl_623 & nor_942_cse;
  assign and_dcpl_1389 = and_dcpl_1383 & and_dcpl_1351 & and_dcpl_1278;
  assign and_dcpl_1391 = and_dcpl_1383 & and_dcpl_73 & and_dcpl_1278;
  assign and_dcpl_1393 = and_dcpl_1349 & and_dcpl_623 & and_dcpl_50;
  assign and_dcpl_1395 = and_dcpl_1383 & and_817_cse & and_dcpl_1278;
  assign and_dcpl_1396 = (~ (fsm_output[7])) & (fsm_output[5]);
  assign and_dcpl_1398 = not_tmp_682 & and_dcpl_1396 & (~ (fsm_output[4]));
  assign and_dcpl_1399 = and_dcpl_623 & (fsm_output[3]);
  assign and_dcpl_1401 = and_dcpl_1399 & nor_668_cse & and_dcpl_1278;
  assign and_dcpl_1404 = and_dcpl_1349 & and_dcpl_623 & and_dcpl_171;
  assign and_dcpl_1406 = and_dcpl_1399 & and_dcpl_1351 & and_dcpl_1278;
  assign and_dcpl_1408 = not_tmp_680 & and_dcpl_1396 & and_dcpl_410;
  assign and_dcpl_1410 = and_dcpl_1399 & and_dcpl_73 & and_dcpl_1278;
  assign and_dcpl_1412 = and_dcpl_1399 & and_817_cse & and_dcpl_1278;
  assign nor_409_nl = ~((fsm_output[3:1]!=3'b000) | (~ nor_tmp_216));
  assign nor_410_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[2])) | (~ (fsm_output[3]))
      | (fsm_output[4]) | (fsm_output[6]));
  assign mux_985_nl = MUX_s_1_2_2((nor_409_nl), (nor_410_nl), fsm_output[0]);
  assign and_dcpl_1413 = (mux_985_nl) & and_dcpl_1396;
  assign and_dcpl_1415 = and_dcpl_658 & (~ (fsm_output[3]));
  assign and_dcpl_1417 = and_dcpl_1415 & nor_668_cse & and_dcpl_1278;
  assign and_dcpl_1419 = and_dcpl_1349 & and_dcpl_658 & nor_942_cse;
  assign and_dcpl_1421 = and_dcpl_1415 & and_dcpl_1351 & and_dcpl_1278;
  assign and_dcpl_1423 = not_tmp_680 & and_dcpl_1396 & and_dcpl_1354;
  assign and_dcpl_1425 = and_dcpl_1415 & and_dcpl_73 & and_dcpl_1278;
  assign and_dcpl_1427 = and_dcpl_1349 & and_dcpl_658 & and_dcpl_50;
  assign and_dcpl_1429 = and_dcpl_1415 & and_817_cse & and_dcpl_1278;
  assign and_dcpl_1430 = and_dcpl_658 & (fsm_output[3]);
  assign and_dcpl_1432 = and_dcpl_1430 & nor_668_cse & and_dcpl_1278;
  assign and_dcpl_1434 = and_dcpl_1349 & and_dcpl_658 & and_dcpl_171;
  assign and_dcpl_1436 = and_dcpl_1430 & and_dcpl_1351 & and_dcpl_1278;
  assign and_dcpl_1438 = not_tmp_680 & and_dcpl_1396 & and_862_cse;
  assign and_dcpl_1440 = and_dcpl_1430 & and_dcpl_73 & and_dcpl_1278;
  assign and_dcpl_1442 = and_dcpl_1349 & and_dcpl_658 & and_2650_cse;
  assign and_dcpl_1444 = and_dcpl_1430 & and_817_cse & and_dcpl_1278;
  assign or_1476_nl = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[4])
      | (fsm_output[5]) | (~ (fsm_output[7]));
  assign nand_151_nl = ~((fsm_output[1]) & (fsm_output[2]) & (fsm_output[3]) & (fsm_output[4])
      & (fsm_output[5]) & (~ (fsm_output[7])));
  assign mux_986_nl = MUX_s_1_2_2((or_1476_nl), (nand_151_nl), fsm_output[0]);
  assign and_dcpl_1445 = ~((mux_986_nl) | (fsm_output[6]));
  assign mux_987_nl = MUX_s_1_2_2(or_865_cse_1, or_864_cse, fsm_output[0]);
  assign and_dcpl_1448 = ~((mux_987_nl) | (fsm_output[5]));
  assign and_dcpl_1449 = and_dcpl_1448 & nor_298_cse & nor_668_cse;
  assign and_dcpl_1451 = and_dcpl_1448 & nor_298_cse & and_dcpl_1351;
  assign and_dcpl_1474 = and_dcpl_100 & nor_942_cse & nor_306_cse;
  assign and_dcpl_1476 = and_dcpl_100 & nor_942_cse & and_dcpl_56;
  assign and_dcpl_1483 = and_dcpl_926 & (fsm_output[3:2]==2'b10) & and_dcpl_103;
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_1_or_1_ssc = and_dcpl_1180
      | and_dcpl_1181 | and_dcpl_1184 | and_dcpl_1185 | and_dcpl_1188 | and_dcpl_1190
      | and_dcpl_1192 | and_dcpl_1194 | and_dcpl_1197 | and_dcpl_1199;
  assign nl_SUM_EXP_LOOP_acc_10_sdt = conv_u2u_67_68(CALC_EXP_LOOP_9_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva)
      + conv_u2u_67_68(CALC_EXP_LOOP_10_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva);
  assign SUM_EXP_LOOP_acc_10_sdt = nl_SUM_EXP_LOOP_acc_10_sdt[67:0];
  assign or_tmp_922 = (fsm_output[6]) | (fsm_output[3]) | IndexLoop_stage_0 | (~
      IndexLoop_stage_0_2) | (fsm_output[4]);
  assign not_tmp_1409 = ~((fsm_output[4:3]==2'b11));
  assign not_tmp_1420 = ~((fsm_output[0]) & (fsm_output[2]));
  assign or_tmp_940 = IndexLoop_stage_0 | IndexLoop_stage_0_2;
  assign or_tmp_948 = (fsm_output[7]) | (fsm_output[6]) | (fsm_output[2]) | (~ and_810_cse_1);
  assign or_1621_nl = (fsm_output[2]) | (~ and_810_cse_1);
  assign or_1620_nl = (fsm_output[2:0]!=3'b101);
  assign mux_1093_nl = MUX_s_1_2_2((or_1621_nl), (or_1620_nl), fsm_output[6]);
  assign or_1619_nl = (fsm_output[6]) | nand_210_cse;
  assign mux_1094_nl = MUX_s_1_2_2((mux_1093_nl), (or_1619_nl), fsm_output[7]);
  assign mux_1095_nl = MUX_s_1_2_2((mux_1094_nl), or_tmp_948, IndexLoop_stage_0);
  assign nand_tmp_52 = ~(IndexLoop_stage_0_2 & (~ (mux_1095_nl)));
  assign or_tmp_957 = (fsm_output[7]) | (fsm_output[6]) | (fsm_output[2]) | (~ (fsm_output[1]));
  assign or_1629_nl = (fsm_output[2:1]!=2'b10);
  assign mux_1100_cse = MUX_s_1_2_2(or_1286_cse, (or_1629_nl), fsm_output[6]);
  assign or_1628_nl = (fsm_output[6]) | nand_52_cse;
  assign mux_1101_nl = MUX_s_1_2_2(mux_1100_cse, (or_1628_nl), fsm_output[7]);
  assign mux_1102_nl = MUX_s_1_2_2((mux_1101_nl), or_tmp_957, IndexLoop_stage_0);
  assign nand_tmp_53 = ~(IndexLoop_stage_0_2 & (~ (mux_1102_nl)));
  assign nor_629_nl = ~((fsm_output[2:1]!=2'b01));
  assign nor_630_nl = ~((fsm_output[2:1]!=2'b10));
  assign mux_1134_nl = MUX_s_1_2_2((nor_629_nl), (nor_630_nl), fsm_output[6]);
  assign nor_631_nl = ~((fsm_output[6]) | nand_52_cse);
  assign mux_1135_nl = MUX_s_1_2_2((mux_1134_nl), (nor_631_nl), fsm_output[7]);
  assign nor_632_nl = ~((fsm_output[7]) | (fsm_output[6]) | (fsm_output[2]) | (~
      (fsm_output[1])));
  assign mux_1136_nl = MUX_s_1_2_2((mux_1135_nl), (nor_632_nl), IndexLoop_stage_0);
  assign nand_tmp_54 = ~(IndexLoop_stage_0_2 & (mux_1136_nl));
  assign or_tmp_1095 = (~ (fsm_output[4])) | (fsm_output[6]) | (~ (fsm_output[7]));
  assign or_tmp_1115 = (fsm_output[2]) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[7]);
  assign nor_577_nl = ~(IndexLoop_stage_0 | (fsm_output[2:0]!=3'b101));
  assign mux_1195_nl = MUX_s_1_2_2(nor_649_cse, (nor_577_nl), fsm_output[6]);
  assign nand_tmp_65 = ~(IndexLoop_stage_0_2 & (mux_1195_nl));
  assign or_tmp_1128 = (fsm_output[5]) | (fsm_output[6]) | (fsm_output[2]);
  assign nor_574_nl = ~((fsm_output[5]) | mux_1100_cse);
  assign nor_575_nl = ~((fsm_output[5]) | (fsm_output[6]) | (~ (fsm_output[1])) |
      (fsm_output[2]));
  assign mux_1209_nl = MUX_s_1_2_2((nor_574_nl), (nor_575_nl), IndexLoop_stage_0);
  assign nand_tmp_66 = ~(IndexLoop_stage_0_2 & (mux_1209_nl));
  assign or_tmp_1140 = (fsm_output[6]) | (~ (fsm_output[1])) | (fsm_output[2]);
  assign mux_1214_nl = MUX_s_1_2_2(mux_1100_cse, or_tmp_1140, IndexLoop_stage_0);
  assign nand_tmp_67 = ~(IndexLoop_stage_0_2 & (~ (mux_1214_nl)));
  assign or_1819_nl = (fsm_output[2:0]!=3'b011);
  assign or_1818_nl = (fsm_output[1]) | not_tmp_1420;
  assign mux_tmp_1215 = MUX_s_1_2_2((or_1819_nl), (or_1818_nl), fsm_output[6]);
  assign or_1823_nl = (fsm_output[3]) | mux_tmp_1215;
  assign or_1822_nl = (fsm_output[3]) | (fsm_output[6]) | (~ and_2642_cse);
  assign mux_tmp_1216 = MUX_s_1_2_2((or_1823_nl), (or_1822_nl), fsm_output[7]);
  assign SUM_EXP_LOOP_nor_itm = ~(and_1134_cse | and_dcpl_964);
  assign ReuseLoop_nor_itm = ~(and_1161_cse | and_dcpl_992);
  assign ReuseLoop_mux1h_3_nl = MUX1HOT_s_1_10_2(nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_1_sva_1,
      MultLoop_2_and_5_itm_1, MultLoop_2_and_6_itm_1, MultLoop_2_and_7_itm_1, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_5_sva,
      nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_6_sva, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_7_sva,
      nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_8_sva, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_9_sva,
      nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_sva, {and_1173_cse
      , and_1175_cse , and_1178_cse , and_1180_cse , and_1183_cse , and_1185_cse
      , and_1187_cse , and_1189_cse , and_1193_cse , and_1195_cse});
  assign ReuseLoop_and_2_cse = (ReuseLoop_mux1h_3_nl) & ReuseLoop_nor_itm;
  assign ReuseLoop_or_itm = and_1173_cse | and_1175_cse | and_1178_cse | and_1180_cse
      | and_1183_cse | and_1185_cse | and_1187_cse | and_1189_cse | and_1193_cse
      | and_1195_cse;
  assign IndexLoop_if_nor_itm = ~(and_1173_cse | and_1175_cse | and_1178_cse | and_1180_cse
      | and_1183_cse | and_1185_cse | and_1187_cse | and_1189_cse | and_1193_cse
      | and_1195_cse);
  assign ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_7_cse
      = MUX1HOT_s_1_10_2((~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_1_sva_1),
      (~ MultLoop_2_and_5_itm_1), (~ MultLoop_2_and_6_itm_1), (~ MultLoop_2_and_7_itm_1),
      (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_5_sva), (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_6_sva),
      (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_7_sva), (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_8_sva),
      (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_9_sva), (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_sva),
      {and_1270_cse , and_1273_cse , and_1276_cse , and_1279_cse , and_1282_cse ,
      and_1284_cse , and_1286_cse , and_1288_cse , and_1193_cse , and_1195_cse});
  assign ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_10_cse
      = MUX1HOT_s_1_10_2(nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_1_sva_1,
      MultLoop_2_and_5_itm_1, MultLoop_2_and_6_itm_1, MultLoop_2_and_7_itm_1, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_5_sva,
      nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_6_sva, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_7_sva,
      nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_8_sva, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_9_sva,
      nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_sva, {and_1270_cse
      , and_1273_cse , and_1276_cse , and_1279_cse , and_1282_cse , and_1284_cse
      , and_1286_cse , and_1288_cse , and_1193_cse , and_1195_cse});
  assign ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_2_cse
      = MUX1HOT_s_1_10_2((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg[2]),
      (reg_MultLoop_1_mux_64_itm_1_reg[5]), (reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_reg[5]),
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_1_ftd,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_1_ftd,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_1_ftd,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd,
      (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2[17]),
      {and_1270_cse , and_1273_cse , and_1276_cse , and_1279_cse , and_1282_cse ,
      and_1284_cse , and_1286_cse , and_1288_cse , and_1193_cse , and_1195_cse});
  assign operator_18_8_true_AC_TRN_AC_WRAP_1_or_itm = and_1173_cse | and_1175_cse
      | and_1178_cse | and_1180_cse | and_1183_cse | and_1185_cse | and_1187_cse
      | and_1189_cse | and_dcpl_1474 | and_dcpl_1476;
  assign SUM_EXP_LOOP_nor_2_itm = ~(and_dcpl_1483 | and_1282_cse | and_1193_cse |
      and_1286_cse);
  always @(posedge clk) begin
    if ( rst ) begin
      reg_w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_0_cse <= 1'b0;
      reg_w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_0_cse <= 1'b0;
      reg_w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_0_cse <= 1'b0;
      reg_const_size_out_1_rsci_ivld_core_psct_cse <= 1'b0;
      reg_layer7_out_rsci_ivld_core_psct_cse <= 1'b0;
      InitAccumLoop_1_iacc_6_0_sva_5_0 <= 6'b000000;
      IndexLoop_asn_3_itm_1 <= 1'b0;
      IndexLoop_stage_0 <= 1'b0;
      IndexLoop_stage_0_2 <= 1'b0;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc15_sva
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc0_sva
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc13_sva
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc12_sva
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc11_sva
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc10_sva
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc9_sva
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc8_sva
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc7_sva
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc6_sva
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc5_sva
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc4_sva
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc3_sva
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc2_sva
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc1_sva
          <= 6'b000000;
      InitAccumLoop_2_iacc_3_0_sva <= 4'b0000;
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1
          <= 5'b00000;
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_out_index_3_0_sva_1_2
          <= 1'b0;
      MultLoop_2_MultLoop_2_nor_2_itm_1 <= 1'b0;
      MultLoop_2_and_15_itm_1 <= 1'b0;
      MultLoop_2_and_14_itm_1 <= 1'b0;
      ReuseLoop_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_outidx_const_assign_1_ReuseLoop_2_asn_tmp_3_2_0_psp_sva_1
          <= 3'b000;
      MultLoop_2_and_5_itm_1 <= 1'b0;
      SUM_EXP_LOOP_acc_itm_69_68 <= 2'b00;
    end
    else if ( core_wen ) begin
      reg_w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_0_cse <= and_73_rmff;
      reg_w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_0_cse <= and_dcpl_77;
      reg_w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_0_cse <= and_dcpl_82;
      reg_const_size_out_1_rsci_ivld_core_psct_cse <= ~((mux_471_nl) | or_1398_cse
          | (fsm_output[0]));
      reg_layer7_out_rsci_ivld_core_psct_cse <= and_dcpl_87 & and_817_cse & and_dcpl_94;
      InitAccumLoop_1_iacc_6_0_sva_5_0 <= MUX_v_6_2_2(6'b000000, (InitAccumLoop_1_iacc_mux_nl),
          (nand_149_nl));
      IndexLoop_asn_3_itm_1 <= MUX1HOT_s_1_3_2(IndexLoop_IndexLoop_nor_tmp, (z_out_12[11]),
          (~ z_out_1_3), {and_dcpl_65 , and_dcpl_60 , and_dcpl_55});
      IndexLoop_stage_0 <= (IndexLoop_mux1h_9_nl) | (~((mux_883_nl) | (fsm_output[5])));
      IndexLoop_stage_0_2 <= (~ (mux_688_nl)) & nor_943_cse & (~ (fsm_output[3]))
          & (fsm_output[0]);
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc15_sva
          <= MUX_v_6_2_2(6'b000000, (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_mux_nl),
          and_dcpl_65);
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc0_sva
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc15_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc13_sva
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc12_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc12_sva
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc11_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc11_sva
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc10_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc10_sva
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc9_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc9_sva
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc8_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc8_sva
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc7_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc7_sva
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc6_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc6_sva
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc5_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc5_sva
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc4_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc4_sva
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc3_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc3_sva
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc2_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc2_sva
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc1_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc1_sva
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc0_sva;
      InitAccumLoop_2_iacc_3_0_sva <= MUX_v_4_2_2(4'b0000, z_out_4, (nand_148_nl));
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1
          <= ROM_1i11_1o5_b94ddd86102738ded3ce1c444a799cda31_1;
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_out_index_3_0_sva_1_2
          <= MultLoop_2_1_acc_3_tmp[2];
      MultLoop_2_MultLoop_2_nor_2_itm_1 <= MultLoop_2_and_5_itm;
      MultLoop_2_and_15_itm_1 <= MultLoop_2_and_6_itm;
      MultLoop_2_and_14_itm_1 <= MultLoop_2_and_7_itm;
      ReuseLoop_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_outidx_const_assign_1_ReuseLoop_2_asn_tmp_3_2_0_psp_sva_1
          <= ROM_1i9_1o3_2fa806bf16b3e0d54016201674d036b62f_1;
      MultLoop_2_and_5_itm_1 <= MUX_s_1_2_2(MultLoop_2_and_5_itm, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_2_sva_mx0w1,
          and_dcpl_520);
      SUM_EXP_LOOP_acc_itm_69_68 <= SUM_EXP_LOOP_mux_1_rgt[69:68];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer7_out_rsci_idat_11_0 <= 12'b000000000000;
    end
    else if ( core_wen & ((and_dcpl_87 & and_dcpl_84 & IndexLoop_stage_0 & nnet_softmax_layer6_t_result_t_softmax_config7_for_1_or_tmp)
        | layer7_out_rsci_idat_11_0_mx0c1) ) begin
      layer7_out_rsci_idat_11_0 <= MUX_v_12_2_2(nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_11_0_lpi_2,
          nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000,
          layer7_out_rsci_idat_11_0_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer7_out_rsci_idat_29_18 <= 12'b000000000000;
    end
    else if ( core_wen & ((and_dcpl_101 & and_dcpl_95 & and_dcpl_93) | layer7_out_rsci_idat_29_18_mx0c1)
        ) begin
      layer7_out_rsci_idat_29_18 <= MUX_v_12_2_2(nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000,
          nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_29_18_lpi_2,
          layer7_out_rsci_idat_29_18_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer7_out_rsci_idat_47_36 <= 12'b000000000000;
    end
    else if ( core_wen & ((and_dcpl_101 & and_dcpl_95 & and_dcpl_109 & (~ (InitAccumLoop_2_iacc_3_0_sva[0])))
        | layer7_out_rsci_idat_47_36_mx0c1) ) begin
      layer7_out_rsci_idat_47_36 <= MUX_v_12_2_2(nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000,
          nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_47_36_lpi_2,
          layer7_out_rsci_idat_47_36_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer7_out_rsci_idat_65_54 <= 12'b000000000000;
    end
    else if ( core_wen & ((and_dcpl_101 & and_dcpl_95 & and_dcpl_109 & (InitAccumLoop_2_iacc_3_0_sva[0]))
        | layer7_out_rsci_idat_65_54_mx0c1) ) begin
      layer7_out_rsci_idat_65_54 <= MUX_v_12_2_2(nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000,
          nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_65_54_lpi_2,
          layer7_out_rsci_idat_65_54_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer7_out_rsci_idat_83_72 <= 12'b000000000000;
    end
    else if ( core_wen & ((and_dcpl_101 & and_dcpl_95 & and_dcpl_120 & (~ (InitAccumLoop_2_iacc_3_0_sva[0])))
        | layer7_out_rsci_idat_83_72_mx0c1) ) begin
      layer7_out_rsci_idat_83_72 <= MUX_v_12_2_2(nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000,
          nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_83_72_lpi_2,
          layer7_out_rsci_idat_83_72_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer7_out_rsci_idat_101_90 <= 12'b000000000000;
    end
    else if ( core_wen & ((and_dcpl_101 & and_dcpl_95 & and_dcpl_120 & (InitAccumLoop_2_iacc_3_0_sva[0]))
        | layer7_out_rsci_idat_101_90_mx0c1) ) begin
      layer7_out_rsci_idat_101_90 <= MUX_v_12_2_2(nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000,
          nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_101_90_lpi_2,
          layer7_out_rsci_idat_101_90_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer7_out_rsci_idat_119_108 <= 12'b000000000000;
    end
    else if ( core_wen & ((and_dcpl_101 & and_dcpl_95 & and_dcpl_131 & (~ (InitAccumLoop_2_iacc_3_0_sva[0])))
        | layer7_out_rsci_idat_119_108_mx0c1) ) begin
      layer7_out_rsci_idat_119_108 <= MUX_v_12_2_2(nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000,
          nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_119_108_lpi_2,
          layer7_out_rsci_idat_119_108_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer7_out_rsci_idat_137_126 <= 12'b000000000000;
    end
    else if ( core_wen & ((and_dcpl_101 & and_dcpl_95 & and_dcpl_131 & (InitAccumLoop_2_iacc_3_0_sva[0]))
        | layer7_out_rsci_idat_137_126_mx0c1) ) begin
      layer7_out_rsci_idat_137_126 <= MUX_v_12_2_2(nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000,
          nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_137_126_lpi_2,
          layer7_out_rsci_idat_137_126_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer7_out_rsci_idat_155_144 <= 12'b000000000000;
    end
    else if ( core_wen & ((and_dcpl_101 & and_dcpl_143 & and_dcpl_92 & (~ (InitAccumLoop_2_iacc_3_0_sva[0])))
        | layer7_out_rsci_idat_155_144_mx0c1) ) begin
      layer7_out_rsci_idat_155_144 <= MUX_v_12_2_2(nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000,
          nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_155_144_lpi_2,
          layer7_out_rsci_idat_155_144_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer7_out_rsci_idat_173_162 <= 12'b000000000000;
    end
    else if ( core_wen & ((and_dcpl_101 & and_dcpl_143 & and_dcpl_93) | layer7_out_rsci_idat_173_162_mx0c1)
        ) begin
      layer7_out_rsci_idat_173_162 <= MUX_v_12_2_2(nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000,
          nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_173_162_lpi_2,
          layer7_out_rsci_idat_173_162_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b11110) & core_wen
        & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_1_1_sva_1 <= 18'b000000000000000000;
    end
    else if ( nor_936_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[1:0]==2'b01) & nor_937_cse
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_1_1_sva_1 <= MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_1_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_61_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b11101) & core_wen
        & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_61_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_61_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_sva_1 <= 18'b000000000000000000;
    end
    else if ( nor_936_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[1:0]==2'b10) & nor_937_cse
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_sva_1 <= MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_60_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[2]) & nor_923_cse &
        (InitAccumLoop_1_iacc_6_0_sva_5_0[4:3]==2'b11) & core_wen & (fsm_output[1])
        & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_60_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_60_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_sva_1 <= 18'b000000000000000000;
    end
    else if ( nor_936_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[1:0]==2'b11) & nor_937_cse
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_sva_1 <= MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_59_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b11011) & core_wen
        & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_59_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_59_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_sva_1 <= 18'b000000000000000000;
    end
    else if ( (~ mux_990_cse) & (InitAccumLoop_1_iacc_6_0_sva_5_0[2]) & nor_923_cse
        & nor_937_cse & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse &
        nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_sva_1 <= MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_58_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b11010) & core_wen
        & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_58_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_58_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_sva_1 <= 18'b000000000000000000;
    end
    else if ( (~ mux_990_cse) & (InitAccumLoop_1_iacc_6_0_sva_5_0[2:0]==3'b101) &
        nor_937_cse & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_sva_1 <= MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b11001) & core_wen
        & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_6_1_sva_1 <= 18'b000000000000000000;
    end
    else if ( (~ mux_990_cse) & (InitAccumLoop_1_iacc_6_0_sva_5_0[2:0]==3'b110) &
        nor_937_cse & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_6_1_sva_1 <= MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_6_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[2])) & nor_923_cse
        & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:3]==2'b11) & core_wen & (fsm_output[1])
        & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_sva_1 <= 18'b000000000000000000;
    end
    else if ( (~ mux_990_cse) & (InitAccumLoop_1_iacc_6_0_sva_5_0[2:0]==3'b111) &
        nor_937_cse & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_sva_1 <= MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b10111) & core_wen
        & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_8_1_sva_1 <= 18'b000000000000000000;
    end
    else if ( nor_936_cse & nor_923_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:3]==2'b01)
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_8_1_sva_1 <= MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_8_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b10110) & core_wen
        & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_9_1_sva_1 <= 18'b000000000000000000;
    end
    else if ( nor_936_cse & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[1])) & (InitAccumLoop_1_iacc_6_0_sva_5_0[0])
        & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[4])) & (InitAccumLoop_1_iacc_6_0_sva_5_0[3])
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_9_1_sva_1 <= MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_9_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b10101) & core_wen
        & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_10_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( nor_936_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[1]) & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[0]))
        & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[4])) & (InitAccumLoop_1_iacc_6_0_sva_5_0[3])
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_10_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_10_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[2]) & nor_923_cse &
        (InitAccumLoop_1_iacc_6_0_sva_5_0[4:3]==2'b10) & core_wen & (fsm_output[1])
        & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( nor_936_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[1]) & (InitAccumLoop_1_iacc_6_0_sva_5_0[0])
        & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[4])) & (InitAccumLoop_1_iacc_6_0_sva_5_0[3])
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b10011) & core_wen
        & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( (~ mux_990_cse) & (InitAccumLoop_1_iacc_6_0_sva_5_0[2]) & nor_923_cse
        & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:3]==2'b01) & core_wen & (fsm_output[1])
        & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b10010) & core_wen
        & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( (~ mux_990_cse) & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b01101)
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b10001) & core_wen
        & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( (~ mux_990_cse) & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b01110)
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[2])) & nor_923_cse
        & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:3]==2'b10) & core_wen & (fsm_output[1])
        & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( (~ mux_990_cse) & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b01111)
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b01111) & core_wen
        & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( nor_936_cse & nor_923_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:3]==2'b10)
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b01110) & core_wen
        & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( nor_936_cse & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[1])) & (InitAccumLoop_1_iacc_6_0_sva_5_0[0])
        & (InitAccumLoop_1_iacc_6_0_sva_5_0[4]) & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[3]))
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b01101) & core_wen
        & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( nor_936_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[1]) & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[0]))
        & (InitAccumLoop_1_iacc_6_0_sva_5_0[4]) & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[3]))
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[2]) & nor_923_cse &
        (InitAccumLoop_1_iacc_6_0_sva_5_0[4:3]==2'b01) & core_wen & (fsm_output[1])
        & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( nor_936_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[1]) & (InitAccumLoop_1_iacc_6_0_sva_5_0[0])
        & (InitAccumLoop_1_iacc_6_0_sva_5_0[4]) & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[3]))
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b01011) & core_wen
        & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( (~ mux_990_cse) & (InitAccumLoop_1_iacc_6_0_sva_5_0[2]) & nor_923_cse
        & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:3]==2'b10) & core_wen & (fsm_output[1])
        & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b01010) & core_wen
        & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( (~ mux_990_cse) & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b10101)
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b01001) & core_wen
        & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( (~ mux_990_cse) & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b10110)
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[2])) & nor_923_cse
        & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:3]==2'b01) & core_wen & (fsm_output[1])
        & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( (~ mux_990_cse) & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b10111)
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[2:0]==3'b111) & nor_937_cse
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( nor_936_cse & nor_923_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:3]==2'b11)
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[2:0]==3'b110) & nor_937_cse
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( nor_936_cse & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[1])) & (InitAccumLoop_1_iacc_6_0_sva_5_0[0])
        & (InitAccumLoop_1_iacc_6_0_sva_5_0[4]) & (InitAccumLoop_1_iacc_6_0_sva_5_0[3])
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[2:0]==3'b101) & nor_937_cse
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( nor_936_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[1]) & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[0]))
        & (InitAccumLoop_1_iacc_6_0_sva_5_0[4]) & (InitAccumLoop_1_iacc_6_0_sva_5_0[3])
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[2]) & nor_923_cse &
        nor_937_cse & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( nor_936_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[1]) & (InitAccumLoop_1_iacc_6_0_sva_5_0[0])
        & (InitAccumLoop_1_iacc_6_0_sva_5_0[4]) & (InitAccumLoop_1_iacc_6_0_sva_5_0[3])
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[2:0]==3'b011) & nor_937_cse
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( (~ mux_990_cse) & (InitAccumLoop_1_iacc_6_0_sva_5_0[2]) & nor_923_cse
        & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:3]==2'b11) & core_wen & (fsm_output[1])
        & nor_942_cse & nor_943_cse & nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[2:0]==3'b010) & nor_937_cse
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( (~ mux_990_cse) & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b11101)
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (InitAccumLoop_1_iacc_6_0_sva_5_0[2:0]==3'b001) & nor_937_cse
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( (~ mux_990_cse) & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b11110)
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( mux_989_cse & (~ (InitAccumLoop_1_iacc_6_0_sva_5_0[2])) & nor_923_cse
        & nor_937_cse & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse &
        nor_944_cse ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_sva_1 <=
          18'b000000000000000000;
    end
    else if ( (~ mux_990_cse) & (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]==5'b11111)
        & core_wen & (fsm_output[1]) & nor_942_cse & nor_943_cse & nor_944_cse )
        begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_sva_1 <=
          MUX_v_18_2_2(InitAccumLoop_slc_InitAccumLoop_iacc_slc_InitAccumLoop_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_sva_1_mx2,
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_62_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_366 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_385_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_62_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_385_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_61_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_377 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_383_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_61_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_383_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_60_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_383 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_381_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_60_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_381_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_59_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_386 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_379_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_59_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_379_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_58_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_389 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_377_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_58_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_377_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_57_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_392 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_375_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_57_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_375_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_56_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_395 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_373_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_56_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_373_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_55_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_398 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_371_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_55_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_371_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_54_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_402 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_369_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_54_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_369_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_53_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_405 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_367_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_53_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_367_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_52_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_407 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_365_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_52_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_365_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_51_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_409 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_363_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_51_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_363_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_50_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_411 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_361_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_50_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_361_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_49_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_413 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_359_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_49_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_359_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_48_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_415 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_357_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_48_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_357_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_47_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_417 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_355_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_47_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_355_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_46_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_419 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_353_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_46_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_353_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_45_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_421 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_351_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_45_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_351_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_44_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_423 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_349_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_44_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_349_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_43_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_425 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_347_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_43_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_347_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_42_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_427 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_345_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_42_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_345_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_41_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_429 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_343_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_41_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_343_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_40_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_431 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_341_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_40_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_341_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_39_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_433 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_339_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_39_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_339_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_38_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_435 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_337_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_38_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_337_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_37_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_437 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_335_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_37_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_335_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_36_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_439 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_333_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_36_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_333_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_35_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_441 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_331_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_35_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_331_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_34_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_443 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_329_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_34_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_329_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_33_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_445 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_327_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_33_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_327_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_32_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_447 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_325_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_32_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_325_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_1_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_372 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_327_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_1_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_327_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_2_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_382 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_329_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_2_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_329_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_3_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_384 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_331_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_3_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_331_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_4_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_388 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_333_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_4_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_333_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_5_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_390 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_335_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_5_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_335_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_6_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_394 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_337_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_6_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_337_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_7_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_396 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_339_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_7_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_339_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_8_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_400 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_341_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_8_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_341_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_9_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_404 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_343_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_9_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_343_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_10_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_406 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_345_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_10_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_345_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_11_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_408 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_347_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_11_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_347_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_12_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_410 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_349_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_12_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_349_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_13_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_412 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_351_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_13_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_351_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_14_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_414 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_353_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_14_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_353_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_15_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_416 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_355_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_15_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_355_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_16_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_418 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_357_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_16_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_357_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_17_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_420 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_359_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_17_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_359_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_18_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_422 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_361_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_18_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_361_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_19_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_424 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_363_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_19_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_363_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_20_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_426 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_365_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_20_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_365_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_21_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_428 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_367_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_21_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_367_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_22_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_430 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_369_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_22_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_369_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_23_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_432 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_371_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_23_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_371_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_24_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_434 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_373_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_24_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_373_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_25_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_436 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_375_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_25_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_375_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_26_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_438 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_377_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_26_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_377_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_27_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_440 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_379_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_27_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_379_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_28_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_442 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_381_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_28_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_381_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_29_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_444 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_383_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_29_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_383_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_30_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_446 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_385_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_30_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_385_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_31_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_cse
        & ((~(or_dcpl_448 | and_dcpl_60)) | nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_263_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_31_sva_1 <= MUX_v_18_2_2(InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_263_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_8_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_cse
        & ((~(or_dcpl_351 | and_dcpl_55)) | nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_57_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_8_sva_1 <= MUX_v_18_2_2(InitAccumLoop_2_slc_InitAccumLoop_2_asn_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_57_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_7_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_cse
        & ((~(or_dcpl_349 | and_dcpl_55)) | nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_53_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_7_sva_1 <= MUX_v_18_2_2(InitAccumLoop_2_slc_InitAccumLoop_2_asn_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_53_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_6_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_cse
        & ((~(or_dcpl_348 | and_dcpl_55)) | nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_49_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_6_sva_1 <= MUX_v_18_2_2(InitAccumLoop_2_slc_InitAccumLoop_2_asn_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_49_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_5_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_cse
        & ((~(or_dcpl_347 | and_dcpl_55)) | nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_45_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_5_sva_1 <= MUX_v_18_2_2(InitAccumLoop_2_slc_InitAccumLoop_2_asn_18_17_0_ctmp_sva_1,
          z_out_20, nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_45_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_1_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_cse
        & ((~(or_dcpl_339 | and_dcpl_55)) | nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_41_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_1_sva_1 <= MUX_v_18_2_2(InitAccumLoop_2_slc_InitAccumLoop_2_asn_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_41_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_2_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_cse
        & ((~(or_dcpl_341 | and_dcpl_55)) | nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_37_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_2_sva_1 <= MUX_v_18_2_2(InitAccumLoop_2_slc_InitAccumLoop_2_asn_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_37_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_3_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_cse
        & ((~(or_dcpl_343 | and_dcpl_55)) | nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_33_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_3_sva_1 <= MUX_v_18_2_2(InitAccumLoop_2_slc_InitAccumLoop_2_asn_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_33_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_4_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_cse
        & ((~(or_dcpl_346 | and_dcpl_55)) | nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_29_rgt)
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_4_sva_1 <= MUX_v_18_2_2(InitAccumLoop_2_slc_InitAccumLoop_2_asn_18_17_0_ctmp_sva_1,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_and_29_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc1_sva_1
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc2_sva_1
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc3_sva_1
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc4_sva_1
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc5_sva_1
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc6_sva_1
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc7_sva_1
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc8_sva_1
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc9_sva_1
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc10_sva_1
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc11_sva_1
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc12_sva_1
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc13_sva_1
          <= 6'b000000;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc14_sva_1
          <= 6'b000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_and_cse
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc1_sva_1
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc0_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc2_sva_1
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc1_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc3_sva_1
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc2_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc4_sva_1
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc3_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc5_sva_1
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc4_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc6_sva_1
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc5_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc7_sva_1
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc6_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc8_sva_1
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc7_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc9_sva_1
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc8_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc10_sva_1
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc9_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc11_sva_1
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc10_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc12_sva_1
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc11_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc13_sva_1
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc12_sva;
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc14_sva_1
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc13_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_101_90_lpi_2
          <= 12'b000000000000;
    end
    else if ( nnet_softmax_layer6_t_result_t_softmax_config7_for_1_and_cse & (~(or_dcpl_472
        | or_dcpl_337)) ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_101_90_lpi_2
          <= nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_119_108_lpi_2
          <= 12'b000000000000;
    end
    else if ( nnet_softmax_layer6_t_result_t_softmax_config7_for_1_and_cse & (~(or_dcpl_472
        | or_dcpl_340)) ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_119_108_lpi_2
          <= nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_11_0_lpi_2
          <= 12'b000000000000;
    end
    else if ( core_wen & (~(or_dcpl_334 | (fsm_output[4:3]!=2'b11) | nand_52_cse
        | (fsm_output[0]) | (~ IndexLoop_stage_0) | nnet_softmax_layer6_t_result_t_softmax_config7_for_1_or_tmp))
        ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_11_0_lpi_2
          <= nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_137_126_lpi_2
          <= 12'b000000000000;
    end
    else if ( nnet_softmax_layer6_t_result_t_softmax_config7_for_1_and_cse & (~(or_dcpl_472
        | or_dcpl_342)) ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_137_126_lpi_2
          <= nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_155_144_lpi_2
          <= 12'b000000000000;
    end
    else if ( nnet_softmax_layer6_t_result_t_softmax_config7_for_1_and_cse & (~(or_dcpl_481
        | or_dcpl_344)) ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_155_144_lpi_2
          <= nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_173_162_lpi_2
          <= 12'b000000000000;
    end
    else if ( nnet_softmax_layer6_t_result_t_softmax_config7_for_1_and_cse & (~(or_dcpl_481
        | or_dcpl_337)) ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_173_162_lpi_2
          <= nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_29_18_lpi_2
          <= 12'b000000000000;
    end
    else if ( nnet_softmax_layer6_t_result_t_softmax_config7_for_1_and_cse & (~(or_dcpl_484
        | or_dcpl_337)) ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_29_18_lpi_2
          <= nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_47_36_lpi_2
          <= 12'b000000000000;
    end
    else if ( nnet_softmax_layer6_t_result_t_softmax_config7_for_1_and_cse & (~(or_dcpl_484
        | or_dcpl_340)) ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_47_36_lpi_2
          <= nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_65_54_lpi_2
          <= 12'b000000000000;
    end
    else if ( nnet_softmax_layer6_t_result_t_softmax_config7_for_1_and_cse & (~(or_dcpl_484
        | or_dcpl_342)) ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_65_54_lpi_2
          <= nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_83_72_lpi_2
          <= 12'b000000000000;
    end
    else if ( nnet_softmax_layer6_t_result_t_softmax_config7_for_1_and_cse & (~(or_dcpl_472
        | or_dcpl_344)) ) begin
      nnet_softmax_layer6_t_result_t_softmax_config7_for_1_io_read_layer7_out_rsc_sdt_83_72_lpi_2
          <= nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_res_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_slc_nnet_softmax_layer6_t_result_t_softmax_config7_for_1_i_3_0_tmp_1000000;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg <=
          3'b000;
    end
    else if ( (mux_1057_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg <=
          nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_192_rgt[17:15];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_1_reg
          <= 3'b000;
    end
    else if ( (mux_1064_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_1_reg
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_192_rgt[14:12];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_2_reg
          <= 12'b000000000000;
    end
    else if ( (mux_1071_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_2_reg
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_192_rgt[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_63_1_ftd <=
          1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_63_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_63_1_ftd <=
          MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (reg_MultLoop_1_mux_64_itm_1_reg[5]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_8_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_272_rgt
          , MultLoop_and_251_rgt , MultLoop_and_252_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_642_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_63_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_63_ssc
        & ((mux_934_nl) | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_491_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_63_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), ({(reg_MultLoop_1_mux_64_itm_1_reg[4:0])
          , reg_MultLoop_1_mux_64_itm_1_1_reg}), (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_8_sva_1[16:0]),
          ({nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12
          , nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0}),
          ({nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12
          , nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0}),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_272_rgt
          , MultLoop_and_251_rgt , MultLoop_and_252_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_642_rgt
          , (and_591_nl) , (and_593_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_64_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_7_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_271_rgt
          , MultLoop_and_243_rgt , MultLoop_and_244_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_637_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_64_ssc
        & (~((~ mux_tmp_500) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_482_m1c))
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_7_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_16_0_lpi_1_dfm_mx0w2,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_271_rgt
          , MultLoop_and_243_rgt , MultLoop_and_244_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_637_rgt
          , (and_587_nl) , (and_588_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_61_1_sva_2 <=
          18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_65_cse
        & (and_225_rgt | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_304_rgt
        | MultLoop_and_242_rgt | and_232_rgt) ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_61_1_sva_2 <=
          MUX1HOT_v_18_4_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_61_1_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_62_sva_1,
          {and_225_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_304_rgt
          , MultLoop_and_242_rgt , and_232_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_65 | and_dcpl_60 | (~ (mux_523_nl)) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_sva_2_mx0c3)
        & (~ nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_243_rgt)
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_20_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_270_rgt
          , MultLoop_and_239_rgt , MultLoop_and_240_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_630_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_16_15
          <= 2'b00;
    end
    else if ( (mux_1074_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_16_15
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_796_rgt[16:15];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_14_0
          <= 15'b000000000000000;
    end
    else if ( (mux_1077_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_14_0
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_796_rgt[14:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_60_1_sva_2 <=
          18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_65_cse
        & (and_243_rgt | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_303_rgt
        | MultLoop_and_238_rgt | and_246_rgt) ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_60_1_sva_2 <=
          MUX1HOT_v_18_4_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_60_1_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_61_sva_1,
          {and_243_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_303_rgt
          , MultLoop_and_238_rgt , and_246_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_68_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_30_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_269_rgt
          , MultLoop_and_235_rgt , MultLoop_and_236_rgt , and_254_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_68_ssc
        & (mux_tmp_861 | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_533_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_30_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_269_rgt
          , MultLoop_and_235_rgt , MultLoop_and_236_rgt , and_254_rgt , (and_638_nl)
          , (and_639_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_59_1_sva_2 <=
          18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_65_cse
        & (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_268_rgt
        | MultLoop_and_233_rgt | MultLoop_and_234_rgt | and_261_rgt) ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_59_1_sva_2 <=
          MUX1HOT_v_18_4_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_59_1_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_6_sva_1,
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_268_rgt
          , MultLoop_and_233_rgt , MultLoop_and_234_rgt , and_261_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_70_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_40_sva_1[17]),
          {and_265_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_302_rgt
          , MultLoop_and_232_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_642_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_70_ssc
        & ((mux_950_nl) | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_544_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_40_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_265_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_302_rgt
          , MultLoop_and_232_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_642_rgt
          , (and_662_nl) , (and_664_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_58_1_sva_2 <=
          18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_65_cse
        & (and_268_rgt | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_301_rgt
        | MultLoop_and_230_rgt | and_274_rgt) ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_58_1_sva_2 <=
          MUX1HOT_v_18_4_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_58_1_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_59_sva_1,
          {and_268_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_301_rgt
          , MultLoop_and_230_rgt , and_274_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_72_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_50_sva_1[17]),
          {and_276_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_300_rgt
          , MultLoop_and_228_rgt , and_280_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_72_ssc
        & (mux_tmp_555 | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_556_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_50_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_276_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_300_rgt
          , MultLoop_and_228_rgt , and_280_rgt , (and_685_nl) , (and_686_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_73_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_58_sva_1[17]),
          {and_282_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_299_rgt
          , MultLoop_and_226_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_608_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_73_ssc
        & (~((fsm_output[2]) & (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_sva_2_mx0c2)))
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_58_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_16_0_lpi_1_dfm_mx0w2,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_282_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_299_rgt
          , MultLoop_and_226_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_608_rgt
          , (and_705_nl) , (and_709_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_6_1_sva_2 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_65_cse
        & (and_287_rgt | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_298_rgt
        | MultLoop_and_224_rgt | and_292_rgt) ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_6_1_sva_2 <= MUX1HOT_v_18_4_2(z_out_20,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_6_1_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_60_sva_1,
          {and_287_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_298_rgt
          , MultLoop_and_224_rgt , and_292_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_75_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_57_sva_1[17]),
          {and_294_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_297_rgt
          , MultLoop_and_222_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_601_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_75_ssc
        & ((mux_959_nl) | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_sva_2_mx0c2)))
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_57_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_294_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_297_rgt
          , MultLoop_and_222_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_601_rgt
          , (and_702_nl) , (and_704_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_76_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_9_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_267_rgt
          , MultLoop_and_219_rgt , MultLoop_and_220_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_596_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_76_ssc
        & (mux_tmp_933 | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_571_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_9_sva_1[16:0]),
          ({nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12
          , nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_10
          , nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_9_0}),
          ({nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12
          , nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0}),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_267_rgt
          , MultLoop_and_219_rgt , MultLoop_and_220_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_596_rgt
          , (and_595_nl) , (and_596_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_77_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_56_sva_1[17]),
          {and_305_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_296_rgt
          , MultLoop_and_218_rgt , and_308_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_77_ssc
        & (mux_tmp_419 | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_sva_2_mx0c2)))
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_56_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_16_0_lpi_1_dfm_mx0w2,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_305_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_296_rgt
          , MultLoop_and_218_rgt , and_308_rgt , (and_699_nl) , (and_701_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_78_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_55_sva_1[17]),
          {and_311_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_295_rgt
          , MultLoop_and_214_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_587_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_78_ssc
        & ((mux_958_nl) | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_sva_2_mx0c2)))
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_55_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_311_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_295_rgt
          , MultLoop_and_214_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_587_rgt
          , (and_696_nl) , (and_698_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_79_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_54_sva_1[17]),
          {and_316_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_294_rgt
          , MultLoop_and_210_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_582_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_79_ssc
        & (~(and_dcpl_169 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_472_m1c))
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_54_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_316_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_294_rgt
          , MultLoop_and_210_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_582_rgt
          , (and_693_nl) , (and_695_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_80_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_53_sva_1[17]),
          {and_320_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_293_rgt
          , MultLoop_and_208_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_577_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_80_ssc
        & ((mux_957_nl) | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_595_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_53_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_320_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_293_rgt
          , MultLoop_and_208_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_577_rgt
          , (and_691_nl) , (and_692_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_155 | and_dcpl_65 | (~ (mux_607_nl)) | and_dcpl_60
        | and_dcpl_55 | and_dcpl_324) & (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_567_cse
        | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_640_cse
        | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_569_cse))
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd
          <= MUX1HOT_s_1_5_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_12_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_3_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_266_rgt
          , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_307_rgt
          , MultLoop_and_206_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_571_rgt
          , and_334_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_2_reg
          <= 5'b00000;
    end
    else if ( (~ (mux_1082_nl)) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_2_reg
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_745_rgt[6:2];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_4_reg
          <= 2'b00;
    end
    else if ( (mux_1087_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_4_reg
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_745_rgt[1:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd_2
          <= 10'b0000000000;
    end
    else if ( (mux_1091_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd_2
          <= MUX1HOT_v_10_9_2((ReuseLoop_ReuseLoop_and_nl), (z_out_20[9:0]), (z_out_21[9:0]),
          (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_sva_1[9:0]),
          (nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0[9:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_9_0,
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_12_sva_1[9:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_3_sva_1[9:0]),
          (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_conc_231_itm_11_0[9:0]),
          {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_470_nl)
          , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_266_rgt
          , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_307_rgt
          , MultLoop_and_206_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_946_rgt
          , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_948_rgt
          , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_571_rgt
          , and_334_rgt , and_dcpl_324});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_82_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_52_sva_1[17]),
          {and_336_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_292_rgt
          , MultLoop_and_204_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_630_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_82_ssc
        & (mux_tmp_594 | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_616_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_52_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_336_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_292_rgt
          , MultLoop_and_204_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_630_rgt
          , (and_689_nl) , (and_690_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_1_ftd
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_65 | (~ (mux_623_nl)) | and_dcpl_60 | and_dcpl_55
        | and_dcpl_338) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_136_cse
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_1_ftd
          <= MUX1HOT_s_1_5_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_13_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_4_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_265_rgt
          , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_306_rgt
          , MultLoop_and_202_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_558_rgt
          , and_347_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_2_reg
          <= 5'b00000;
    end
    else if ( (~ (mux_1099_nl)) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_2_reg
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_747_rgt[16:12];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_3_reg
          <= 12'b000000000000;
    end
    else if ( (~ (mux_1106_nl)) & (fsm_output[0]) & (~ (fsm_output[5])) & core_wen
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_3_reg
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_747_rgt[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_84_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_51_sva_1[17]),
          {and_349_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_291_rgt
          , MultLoop_and_200_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_552_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_84_ssc
        & ((mux_956_nl) | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_631_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_51_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_349_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_291_rgt
          , MultLoop_and_200_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_552_rgt
          , (and_687_nl) , (and_688_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_1_ftd
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_65 | (~ (mux_636_nl)) | and_dcpl_60 | and_dcpl_55
        | and_dcpl_353) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_136_cse
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_1_ftd
          <= MUX1HOT_s_1_5_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_14_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_5_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_264_rgt
          , MultLoop_and_197_rgt , MultLoop_and_198_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_546_rgt
          , and_363_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_2_reg
          <= 5'b00000;
    end
    else if ( (mux_1112_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_2_reg
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_748_rgt[16:12];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_3_reg
          <= 12'b000000000000;
    end
    else if ( (mux_1118_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_3_reg
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_748_rgt[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_86_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_5_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_263_rgt
          , MultLoop_and_195_rgt , MultLoop_and_196_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_540_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_86_ssc
        & ((mux_955_nl) | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_643_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_5_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_263_rgt
          , MultLoop_and_195_rgt , MultLoop_and_196_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_540_rgt
          , (and_683_nl) , (and_684_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_1_ftd
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_65 | (~ (mux_647_nl)) | and_dcpl_60 | and_dcpl_55
        | and_dcpl_369) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_136_cse
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_1_ftd
          <= MUX1HOT_s_1_5_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_15_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_6_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_262_rgt
          , MultLoop_and_193_rgt , MultLoop_and_194_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_534_rgt
          , and_376_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_2_reg
          <= 5'b00000;
    end
    else if ( (mux_1124_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_2_reg
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_749_rgt[16:12];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_3_reg
          <= 12'b000000000000;
    end
    else if ( (mux_1129_nl) & (~ (fsm_output[5])) & (fsm_output[0]) & core_wen )
        begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_3_reg
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_749_rgt[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_88_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_49_sva_1[17]),
          {and_377_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_290_rgt
          , MultLoop_and_192_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_528_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_88_ssc
        & (mux_tmp_642 | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_654_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_49_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_377_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_290_rgt
          , MultLoop_and_192_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_528_rgt
          , (and_681_nl) , (and_682_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_65 | (~ (mux_658_nl)) | and_dcpl_60 | and_dcpl_55)
        & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_136_cse
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd
          <= MUX1HOT_s_1_5_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_16_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_7_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_261_rgt
          , MultLoop_and_189_rgt , MultLoop_and_190_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_522_rgt
          , and_387_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( (mux_1133_nl) & nor_959_cse & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd_1
          <= MUX1HOT_v_17_7_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_16_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_7_sva_1[16:0]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_261_rgt
          , MultLoop_and_189_rgt , MultLoop_and_190_rgt , (and_605_nl) , (and_606_nl)
          , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_522_rgt
          , and_387_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_90_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_48_sva_1[17]),
          {and_388_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_289_rgt
          , MultLoop_and_188_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_522_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_90_ssc
        & ((mux_954_nl) | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_665_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_48_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_388_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_289_rgt
          , MultLoop_and_188_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_522_rgt
          , (and_679_nl) , (and_680_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_65 | (~ (mux_671_nl)) | and_dcpl_60 | and_dcpl_55)
        & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_136_cse
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd
          <= MUX1HOT_s_1_5_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_17_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_8_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_260_rgt
          , MultLoop_and_185_rgt , MultLoop_and_186_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_528_rgt
          , and_393_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( (~ (mux_1139_nl)) & (fsm_output[0]) & (~ (fsm_output[5])) & (~ (fsm_output[3]))
        & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd_1
          <= MUX1HOT_v_17_7_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_17_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_acc_8_sva_1[16:0]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_260_rgt
          , MultLoop_and_185_rgt , MultLoop_and_186_rgt , (and_607_nl) , (and_608_nl)
          , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_528_rgt
          , and_393_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_92_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_47_sva_1[17]),
          {and_394_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_288_rgt
          , MultLoop_and_184_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_534_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_92_ssc
        & (mux_tmp_680 | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_681_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_47_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_16_0_lpi_1_dfm_mx0w2,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_394_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_288_rgt
          , MultLoop_and_184_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_534_rgt
          , (and_677_nl) , (and_678_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2 <=
          18'b000000000000000000;
    end
    else if ( core_wen & (and_dcpl_65 | and_dcpl_60 | and_dcpl_160 | and_dcpl_55)
        & (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_639_cse
        | ((~ IndexLoop_stage_0_2) & and_dcpl_60) | (or_1084_tmp & and_dcpl_55)))
        ) begin
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2 <=
          MUX1HOT_v_18_5_2(z_out_20, z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_1,
          nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_18_sva_1,
          InitAccumLoop_2_slc_InitAccumLoop_2_asn_18_17_0_ctmp_sva_1, {(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_259_nl)
          , (MultLoop_and_181_nl) , (MultLoop_and_182_nl) , (and_400_nl) , and_dcpl_160});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_94_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_46_sva_1[17]),
          {and_403_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_287_rgt
          , MultLoop_and_180_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_546_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_94_ssc
        & ((mux_953_nl) | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_692_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_46_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_403_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_287_rgt
          , MultLoop_and_180_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_546_rgt
          , (and_675_nl) , (and_676_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_65 | and_dcpl_60 | (~ (mux_698_nl)) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_sva_2_mx0c3)
        & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_19_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_258_rgt
          , MultLoop_and_177_rgt , MultLoop_and_178_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_552_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_16_15
          <= 2'b00;
    end
    else if ( (mux_1144_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_16_15
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_778_rgt[16:15];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_14_0
          <= 15'b000000000000000;
    end
    else if ( (mux_1147_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_14_0
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_778_rgt[14:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_96_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_45_sva_1[17]),
          {and_409_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_286_rgt
          , MultLoop_and_176_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_558_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_96_ssc
        & (mux_tmp_691 | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_703_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_45_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_409_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_286_rgt
          , MultLoop_and_176_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_558_rgt
          , (and_673_nl) , (and_674_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_65 | and_dcpl_60 | (~ (mux_708_nl)) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_sva_2_mx0c3)
        & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_2_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_257_rgt
          , MultLoop_and_173_rgt , MultLoop_and_174_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_480_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_16_15
          <= 2'b00;
    end
    else if ( (mux_1150_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_16_15
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_776_rgt[16:15];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_14_0
          <= 15'b000000000000000;
    end
    else if ( (mux_1153_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_14_0
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_776_rgt[14:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_98_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_44_sva_1[17]),
          {and_419_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_285_rgt
          , MultLoop_and_172_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_571_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_98_ssc
        & ((mux_952_nl) | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_714_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_44_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_419_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_285_rgt
          , MultLoop_and_172_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_571_rgt
          , (and_671_nl) , (and_672_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_65 | and_dcpl_60 | (~ (mux_717_nl)) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_sva_2_mx0c3)
        & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_21_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_256_rgt
          , MultLoop_and_169_rgt , MultLoop_and_170_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_577_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_16_15
          <= 2'b00;
    end
    else if ( (mux_1157_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_16_15
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_774_rgt[16:15];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_14_0
          <= 15'b000000000000000;
    end
    else if ( (mux_1160_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_14_0
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_774_rgt[14:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_100_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_43_sva_1[17]),
          {and_426_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_284_rgt
          , MultLoop_and_168_rgt , and_430_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_100_ssc
        & (mux_tmp_724 | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_725_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_43_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_426_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_284_rgt
          , MultLoop_and_168_rgt , and_430_rgt , (and_669_nl) , (and_670_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_65 | and_dcpl_60 | (~ (mux_729_nl)) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_sva_2_mx0c3)
        & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_22_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_255_rgt
          , MultLoop_and_165_rgt , MultLoop_and_166_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_582_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_16_15
          <= 2'b00;
    end
    else if ( (mux_1163_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_16_15
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_772_rgt[16:15];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_14_0
          <= 15'b000000000000000;
    end
    else if ( (mux_1166_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_14_0
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_772_rgt[14:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_102_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_42_sva_1[17]),
          {and_435_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_283_rgt
          , MultLoop_and_164_rgt , and_438_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_102_ssc
        & ((mux_951_nl) | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_739_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_42_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_435_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_283_rgt
          , MultLoop_and_164_rgt , and_438_rgt , (and_667_nl) , (and_668_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_65 | and_dcpl_60 | (~ (mux_745_nl)) | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_sva_2_mx0c3)
        & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_23_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_254_rgt
          , MultLoop_and_161_rgt , MultLoop_and_162_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_587_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_16_15
          <= 2'b00;
    end
    else if ( (mux_1169_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_16_15
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_770_rgt[16:15];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_14_0
          <= 15'b000000000000000;
    end
    else if ( (mux_1173_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_14_0
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_770_rgt[14:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_104_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_41_sva_1[17]),
          {and_442_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_282_rgt
          , MultLoop_and_160_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_596_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_104_ssc
        & (mux_tmp_738 | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_753_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_41_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_442_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_282_rgt
          , MultLoop_and_160_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_596_rgt
          , (and_665_nl) , (and_666_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_1_ftd
          <= 3'b000;
    end
    else if ( core_wen & (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_2_mx0c0
        | and_dcpl_65 | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_591_cse
        | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_2_mx0c3
        | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_2_mx0c4
        | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_2_mx0c5)
        & (~ nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_567_cse)
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_1_ftd
          <= MUX1HOT_v_3_5_2((z_out_20[17:15]), (z_out_21[17:15]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_1[17:15]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_24_sva_1[17:15]),
          ({1'b0 , (MultLoop_1_1_MultLoop_1_mux_nl)}), {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_253_rgt
          , MultLoop_and_157_rgt , MultLoop_and_158_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_2_mx0c3
          , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_2_mx0c4});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_2_reg
          <= 3'b000;
    end
    else if ( (~ (mux_1181_nl)) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_2_reg
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_799_rgt[14:12];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg
          <= 12'b000000000000;
    end
    else if ( (mux_1186_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_799_rgt[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_106_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_4_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_252_rgt
          , MultLoop_and_155_rgt , MultLoop_and_156_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_440_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_106_ssc
        & (~((~ mux_tmp_774) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_447_m1c))
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_4_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_252_rgt
          , MultLoop_and_155_rgt , MultLoop_and_156_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_440_rgt
          , (and_658_nl) , (and_659_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd
          <= 3'b000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_107_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd
          <= MUX1HOT_v_3_4_2((z_out_20[17:15]), (z_out_21[17:15]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_1[17:15]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_25_sva_1[17:15]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_251_rgt
          , MultLoop_and_153_rgt , MultLoop_and_154_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_601_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_2_reg
          <= 3'b000;
    end
    else if ( (~ (mux_1191_nl)) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_2_reg
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_766_rgt[3:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_4_reg
          <= 1'b0;
    end
    else if ( (mux_1194_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_4_reg
          <= nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_mux1h_766_rgt[0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2
          <= 11'b00000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_107_ssc
        & (~ and_dcpl_175) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2
          <= MUX1HOT_v_11_8_2((nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_3_14_0[10:0]),
          (z_out_20[10:0]), (z_out_21[10:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_1[10:0]),
          (ReuseLoop_1_ir_ReuseLoop_1_ir_and_nl), (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_25_sva_1[10:0]),
          ({2'b00 , (ReuseLoop_2_ir_ReuseLoop_2_ir_and_nl)}), (CALC_SOFTMAX_LOOP_6_or_cse[10:0]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_444_cse
          , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_251_rgt
          , MultLoop_and_153_rgt , MultLoop_and_154_rgt , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_446_nl)
          , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_601_rgt
          , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_2_mx0c4
          , (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_845_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_108_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_39_sva_1[17]),
          {and_471_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_281_rgt
          , MultLoop_and_152_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_637_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_108_ssc
        & ((mux_949_nl) | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_788_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_39_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_471_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_281_rgt
          , MultLoop_and_152_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_637_rgt
          , (and_656_nl) , (and_657_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_1_ftd
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_65 | and_dcpl_60 | (~ (mux_796_nl))) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_26_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_250_rgt
          , MultLoop_and_149_rgt , MultLoop_and_150_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_608_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( (~ (mux_1198_nl)) & nor_298_cse & (~ (fsm_output[7])) & core_wen )
        begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_26_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_250_rgt
          , MultLoop_and_149_rgt , MultLoop_and_150_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_608_rgt
          , (and_627_nl) , (and_629_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_110_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_38_sva_1[17]),
          {and_475_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_280_rgt
          , MultLoop_and_148_rgt , and_478_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_110_ssc
        & (mux_tmp_787 | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_802_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_38_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_16_0_lpi_1_dfm_mx0w2,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_475_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_280_rgt
          , MultLoop_and_148_rgt , and_478_rgt , (and_654_nl) , (and_655_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_1_ftd
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_65 | and_dcpl_60 | (~ (mux_807_nl))) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_27_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_249_rgt
          , MultLoop_and_145_rgt , MultLoop_and_146_rgt , and_482_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( (~ (mux_1207_nl)) & nor_952_cse & (fsm_output[0]) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_27_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_249_rgt
          , MultLoop_and_145_rgt , MultLoop_and_146_rgt , and_482_rgt , (and_630_nl)
          , (and_631_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_112_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_37_sva_1[17]),
          {and_483_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_279_rgt
          , MultLoop_and_144_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_540_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_112_ssc
        & ((mux_948_nl) | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_815_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_37_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_483_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_279_rgt
          , MultLoop_and_144_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_540_rgt
          , (and_652_nl) , (and_653_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_1_ftd
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_65 | and_dcpl_60 | (~ (mux_822_nl))) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_28_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_248_rgt
          , MultLoop_and_141_rgt , MultLoop_and_142_rgt , and_489_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( (~ (mux_1212_nl)) & nor_298_cse & (~ (fsm_output[7])) & core_wen )
        begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_28_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_248_rgt
          , MultLoop_and_141_rgt , MultLoop_and_142_rgt , and_489_rgt , (and_632_nl)
          , (and_633_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_114_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_36_sva_1[17]),
          {and_490_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_278_rgt
          , MultLoop_and_140_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_440_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_114_ssc
        & (mux_tmp_831 | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_832_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_36_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_490_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_278_rgt
          , MultLoop_and_140_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_440_rgt
          , (and_650_nl) , (and_651_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_1_ftd
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_65 | and_dcpl_60 | (~ (mux_838_nl))) & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_nor_175_cse
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_29_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_247_rgt
          , MultLoop_and_137_rgt , MultLoop_and_138_rgt , and_495_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( (~ (mux_1217_nl)) & nor_952_cse & (fsm_output[0]) & core_wen ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_29_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_16_0_lpi_1_dfm_mx0w2,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_247_rgt
          , MultLoop_and_137_rgt , MultLoop_and_138_rgt , and_495_rgt , (and_634_nl)
          , (and_635_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_116_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_35_sva_1[17]),
          {and_496_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_277_rgt
          , MultLoop_and_136_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_397_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_116_ssc
        & ((mux_947_nl) | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_846_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_35_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_496_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_277_rgt
          , MultLoop_and_136_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_397_rgt
          , (and_648_nl) , (and_649_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_117_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_3_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_246_rgt
          , MultLoop_and_133_rgt , MultLoop_and_134_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_397_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_117_ssc
        & ((mux_944_nl) | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_850_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_3_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_246_rgt
          , MultLoop_and_133_rgt , MultLoop_and_134_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_397_rgt
          , (and_636_nl) , (and_637_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_118_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_34_sva_1[17]),
          {and_502_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_276_rgt
          , MultLoop_and_132_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_480_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_118_ssc
        & (mux_tmp_845 | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_856_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_34_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_502_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_276_rgt
          , MultLoop_and_132_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_480_rgt
          , (and_646_nl) , (and_647_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_119_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_31_sva_1[17]),
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_245_rgt
          , MultLoop_and_129_rgt , MultLoop_and_130_rgt , and_507_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_119_ssc
        & ((mux_945_nl) | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_862_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_31_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_245_rgt
          , MultLoop_and_129_rgt , MultLoop_and_130_rgt , and_507_rgt , (and_640_nl)
          , (and_641_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_120_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_33_sva_1[17]),
          {and_508_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_275_rgt
          , MultLoop_and_128_rgt , and_512_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_120_ssc
        & ((mux_946_nl) | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_867_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_33_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_508_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_275_rgt
          , MultLoop_and_128_rgt , and_512_rgt , (and_644_nl) , (and_645_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_1_ftd
          <= 1'b0;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_121_ssc
        ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_1_ftd
          <= MUX1HOT_s_1_4_2((z_out_20[17]), (z_out_21[17]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_sva_1[17]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_32_sva_1[17]),
          {and_513_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_274_rgt
          , MultLoop_and_126_rgt , and_516_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_1_ftd_1
          <= 17'b00000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_121_ssc
        & (mux_tmp_870 | (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt
        | (~ mux_872_itm)))) ) begin
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_1_ftd_1
          <= MUX1HOT_v_17_6_2((z_out_20[16:0]), (z_out_21[16:0]), (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_sva_1[16:0]),
          (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_32_sva_1[16:0]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          {and_513_rgt , nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_274_rgt
          , MultLoop_and_126_rgt , and_516_rgt , (and_642_nl) , (and_643_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_reg
          <= 6'b000000;
    end
    else if ( (~ (mux_1223_nl)) & (~ (fsm_output[5])) & core_wen ) begin
      reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_reg
          <= MultLoop_mux1h_60_rgt[17:12];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_1_reg
          <= 12'b000000000000;
    end
    else if ( (mux_1227_nl) & (fsm_output[0]) & (~ (fsm_output[3])) & (~ (fsm_output[5]))
        & core_wen ) begin
      reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_1_reg
          <= MultLoop_mux1h_60_rgt[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MultLoop_1_mux_64_itm_1_reg <= 6'b000000;
    end
    else if ( (mux_1235_nl) & (~ (fsm_output[5])) & core_wen ) begin
      reg_MultLoop_1_mux_64_itm_1_reg <= MultLoop_1_mux1h_65_rgt[17:12];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MultLoop_1_mux_64_itm_1_1_reg <= 12'b000000000000;
    end
    else if ( (mux_1241_nl) & nor_959_cse & core_wen ) begin
      reg_MultLoop_1_mux_64_itm_1_1_reg <= MultLoop_1_mux1h_65_rgt[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_0_sva_1 <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_62_cse
        & (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_639_cse
        | (or_dcpl_490 & and_dcpl_158) | (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_126_tmp
        & and_dcpl_60))) ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_0_sva_1 <= MUX1HOT_v_18_4_2(z_out_20,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_8_1_sva_1,
          InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          {(nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_194_nl)
          , (MultLoop_and_215_nl) , (MultLoop_and_216_nl) , (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_136_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_63_sva <= 18'b000000000000000000;
    end
    else if ( nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_62_cse
        & (~(nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_639_cse
        | (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_127_tmp
        & and_dcpl_60))) ) begin
      nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_63_sva <= MUX1HOT_v_18_4_2(z_out_20,
          z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_9_1_sva_1,
          InitAccumLoop_1_slc_InitAccumLoop_1_iacc_slc_InitAccumLoop_1_iacc_6_0_5_0_1_18_17_0_ctmp_sva_1,
          {(and_555_nl) , (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_195_nl)
          , (MultLoop_and_212_nl) , and_dcpl_158});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer3_out_0_16_0_lpi_1_dfm_16_15 <= 2'b00;
      layer3_out_0_16_0_lpi_1_dfm_14_12 <= 3'b000;
    end
    else if ( and_2617_ssc ) begin
      layer3_out_0_16_0_lpi_1_dfm_16_15 <= MUX_v_2_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_cse_16_15,
          (nnet_relu_layer4_t_layer5_t_relu_config5_for_nnet_relu_layer4_t_layer5_t_relu_config5_for_and_cse[16:15]),
          and_558_ssc);
      layer3_out_0_16_0_lpi_1_dfm_14_12 <= MUX_v_3_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_cse_14_12,
          (nnet_relu_layer4_t_layer5_t_relu_config5_for_nnet_relu_layer4_t_layer5_t_relu_config5_for_and_cse[14:12]),
          and_558_ssc);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer3_out_0_16_0_lpi_1_dfm_11_0 <= 12'b000000000000;
    end
    else if ( mux_1243_cse & (~ (fsm_output[5])) & (fsm_output[1]) & (~ (fsm_output[3]))
        & core_wen ) begin
      layer3_out_0_16_0_lpi_1_dfm_11_0 <= MUX1HOT_v_12_4_2(({2'b00 , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd_2}),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_cse_11_0,
          (nnet_relu_layer4_t_layer5_t_relu_config5_for_nnet_relu_layer4_t_layer5_t_relu_config5_for_and_cse[11:0]),
          CALC_SOFTMAX_LOOP_6_or_cse, {and_dcpl_65 , (and_557_nl) , and_558_ssc ,
          (and_560_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_16_0_lpi_1_dfm <=
          17'b00000000000000000;
    end
    else if ( core_wen & (mux_919_nl) ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_16_0_lpi_1_dfm <=
          MUX_v_17_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_16_0_lpi_1_dfm_mx0w2,
          and_562_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_16_0_lpi_1_dfm <=
          17'b00000000000000000;
    end
    else if ( core_wen & (mux_923_nl) ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_16_0_lpi_1_dfm <=
          MUX_v_17_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_16_0_lpi_1_dfm_mx0w2,
          and_564_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_16_0_lpi_1_dfm_16_12
          <= 5'b00000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_16_0_lpi_1_dfm_11_0
          <= 12'b000000000000;
    end
    else if ( nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_2_ssc ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_16_0_lpi_1_dfm_16_12
          <= MUX_v_5_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_12,
          ({nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_cse_16_15
          , nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_cse_14_12}),
          and_566_rgt);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_16_0_lpi_1_dfm_11_0
          <= MUX_v_12_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11_0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_cse_11_0,
          and_566_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_16_0_lpi_1_dfm_ftd
          <= 2'b00;
      reg_nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_16_0_lpi_1_dfm_ftd_1
          <= 15'b000000000000000;
    end
    else if ( nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_3_ssc ) begin
      reg_nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_16_0_lpi_1_dfm_ftd
          <= MUX_v_2_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_16_0_lpi_1_dfm_mx0w2_16_15,
          and_568_rgt);
      reg_nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_16_0_lpi_1_dfm_ftd_1
          <= MUX_v_15_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_16_0_lpi_1_dfm_mx0w2_14_0,
          and_568_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_16_0_lpi_1_dfm <=
          17'b00000000000000000;
    end
    else if ( core_wen & mux_tmp_926 ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_16_0_lpi_1_dfm <=
          MUX_v_17_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_16_0_lpi_1_dfm_mx0w2,
          and_571_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_16_0_lpi_1_dfm <=
          17'b00000000000000000;
    end
    else if ( core_wen & (mux_929_nl) ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_16_0_lpi_1_dfm <=
          MUX_v_17_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_16_0_lpi_1_dfm_mx0w2,
          and_574_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_16_0_lpi_1_dfm <=
          17'b00000000000000000;
    end
    else if ( core_wen & mux_tmp_928 ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_16_0_lpi_1_dfm <=
          MUX_v_17_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_16_0_lpi_1_dfm_mx0w2,
          and_577_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_16_0_lpi_1_dfm <=
          17'b00000000000000000;
    end
    else if ( core_wen & (mux_931_nl) ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_16_0_lpi_1_dfm <=
          MUX_v_17_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_16_0_lpi_1_dfm_mx0w2,
          and_580_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_16_0_lpi_1_dfm <=
          17'b00000000000000000;
    end
    else if ( core_wen & mux_tmp_930 ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_16_0_lpi_1_dfm <=
          MUX_v_17_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          and_583_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_16_0_lpi_1_dfm <=
          17'b00000000000000000;
    end
    else if ( core_wen & (mux_932_nl) ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_16_0_lpi_1_dfm <=
          MUX_v_17_2_2(nnet_relu_layer4_t_layer5_t_relu_config5_for_nnet_relu_layer4_t_layer5_t_relu_config5_for_and_cse,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          and_585_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_16_0_lpi_1_dfm <=
          17'b00000000000000000;
    end
    else if ( core_wen & (mux_938_nl) ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_16_0_lpi_1_dfm <=
          MUX_v_17_2_2(({nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
          , nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_0}),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          and_610_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_16_0_lpi_1_dfm <=
          17'b00000000000000000;
    end
    else if ( core_wen & (mux_800_nl) ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_16_0_lpi_1_dfm <=
          MUX_v_17_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_16_0_lpi_1_dfm_mx0w0,
          ({nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_16_15
          , nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_14_12
          , nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_11
          , nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_16_0_lpi_1_dfm_mx0w0_10_0}),
          and_624_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MultLoop_2_and_7_itm_1 <= 1'b0;
      MultLoop_2_and_6_itm_1 <= 1'b0;
    end
    else if ( MultLoop_2_and_cse ) begin
      MultLoop_2_and_7_itm_1 <= MUX_s_1_2_2(MultLoop_2_and_7_itm, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_4_sva_mx0w1,
          and_dcpl_520);
      MultLoop_2_and_6_itm_1 <= MUX_s_1_2_2(MultLoop_2_and_6_itm, nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_3_sva_mx0w1,
          and_dcpl_520);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_10_18_6_true_AC_TRN_AC_SAT_18_2_AC_TRN_AC_SAT_exp_arr_0_sva
          <= 67'b0000000000000000000000000000000000000000000000000000000000000000000;
      nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_sva <= 1'b0;
      nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_9_sva <= 1'b0;
      nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_8_sva <= 1'b0;
      nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_7_sva <= 1'b0;
      nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_6_sva <= 1'b0;
      nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_5_sva <= 1'b0;
    end
    else if ( ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_10_18_6_true_AC_TRN_AC_SAT_18_2_AC_TRN_AC_SAT_exp_arr_and_cse
        ) begin
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_10_18_6_true_AC_TRN_AC_SAT_18_2_AC_TRN_AC_SAT_exp_arr_0_sva
          <= z_out_9;
      nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_sva <= nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_sva_mx0w0;
      nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_9_sva <= nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_9_sva_mx0w0;
      nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_8_sva <= nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_8_sva_mx0w0;
      nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_7_sva <= nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_7_sva_mx0w0;
      nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_6_sva <= nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_6_sva_mx0w0;
      nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_5_sva <= nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_5_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CALC_EXP_LOOP_2_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva <= 67'b0000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( core_wen & (~(or_dcpl_455 | or_dcpl_607 | or_dcpl_611)) ) begin
      CALC_EXP_LOOP_2_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva <= z_out_9;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CALC_EXP_LOOP_3_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva <= 67'b0000000000000000000000000000000000000000000000000000000000000000000;
      SUM_EXP_LOOP_acc_9_itm <= 68'b00000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( operator_67_47_false_AC_TRN_AC_WRAP_and_1_cse ) begin
      CALC_EXP_LOOP_3_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva <= z_out_9;
      SUM_EXP_LOOP_acc_9_itm <= z_out_24[67:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CALC_EXP_LOOP_4_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva <= 67'b0000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( core_wen & (~(or_dcpl_455 | or_dcpl_607 | nand_209_cse)) ) begin
      CALC_EXP_LOOP_4_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva <= z_out_9;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CALC_EXP_LOOP_5_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva <= 67'b0000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( core_wen & (~(or_dcpl_455 | or_dcpl_466 | or_1875_cse)) ) begin
      CALC_EXP_LOOP_5_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva <= z_out_9;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      SUM_EXP_LOOP_acc_itm_67_0 <= 68'b00000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ((mux_1247_nl) | (fsm_output[1]) | (~ (fsm_output[0])) | (fsm_output[5])
        | (fsm_output[6]) | (~ (fsm_output[7]))) & core_wen ) begin
      SUM_EXP_LOOP_acc_itm_67_0 <= SUM_EXP_LOOP_mux_1_rgt[67:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CALC_EXP_LOOP_6_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva <= 67'b0000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( core_wen & (~(or_dcpl_455 | or_dcpl_466 | or_dcpl_611)) ) begin
      CALC_EXP_LOOP_6_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva <= z_out_9;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CALC_EXP_LOOP_7_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva <= 67'b0000000000000000000000000000000000000000000000000000000000000000000;
      SUM_EXP_LOOP_acc_11_itm <= 69'b000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( operator_67_47_false_AC_TRN_AC_WRAP_and_5_cse ) begin
      CALC_EXP_LOOP_7_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva <= z_out_9;
      SUM_EXP_LOOP_acc_11_itm <= z_out_10[68:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CALC_EXP_LOOP_8_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva <= 67'b0000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( core_wen & (~(or_dcpl_455 | or_dcpl_466 | nand_209_cse)) ) begin
      CALC_EXP_LOOP_8_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva <= z_out_9;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CALC_EXP_LOOP_9_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva <= 67'b0000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( core_wen & (~(or_dcpl_469 | or_647_cse_1 | or_1875_cse)) ) begin
      CALC_EXP_LOOP_9_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva <= z_out_9;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CALC_EXP_LOOP_10_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva <= 67'b0000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( core_wen & (~(or_dcpl_469 | or_647_cse_1 | or_dcpl_611)) ) begin
      CALC_EXP_LOOP_10_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva <= z_out_9;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_71_51_false_AC_TRN_AC_WRAP_91_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1_dfm
          <= 91'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( core_wen & (~(or_dcpl_469 | or_647_cse_1 | nand_209_cse)) ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_71_51_false_AC_TRN_AC_WRAP_91_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1_dfm
          <= MUX_v_91_2_2(operator_91_21_false_AC_TRN_AC_WRAP_rshift_itm, 91'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
          (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_nor_nl));
    end
  end
  assign or_1411_nl = (fsm_output[2]) | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[7]);
  assign nand_61_nl = ~((fsm_output[2]) & (fsm_output[3]) & (fsm_output[4]) & (fsm_output[7]));
  assign mux_470_nl = MUX_s_1_2_2((or_1411_nl), (nand_61_nl), fsm_output[1]);
  assign or_713_nl = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[4])
      | (fsm_output[7]);
  assign mux_471_nl = MUX_s_1_2_2((mux_470_nl), (or_713_nl), IndexLoop_stage_0);
  assign InitAccumLoop_1_iacc_mux_nl = MUX_v_6_2_2((z_out[5:0]), IndexLoop_mux_1_tmp,
      and_dcpl_65);
  assign nand_99_nl = ~((fsm_output[1]) & (fsm_output[2]) & (~ (fsm_output[6])) &
      (fsm_output[7]));
  assign mux_152_nl = MUX_s_1_2_2(or_381_cse, or_1298_cse, fsm_output[1]);
  assign mux_477_nl = MUX_s_1_2_2((nand_99_nl), (mux_152_nl), z_out[6]);
  assign or_378_nl = (fsm_output[2]) | (fsm_output[6]) | (fsm_output[7]);
  assign or_377_nl = (fsm_output[2]) | (~ (fsm_output[6])) | (fsm_output[7]);
  assign mux_151_nl = MUX_s_1_2_2((or_378_nl), (or_377_nl), fsm_output[1]);
  assign mux_478_nl = MUX_s_1_2_2((mux_477_nl), (mux_151_nl), fsm_output[0]);
  assign nand_149_nl = ~((~ (mux_478_nl)) & and_dcpl_169);
  assign nnet_dense_large_input_t_layer2_t_config2_if_nnet_dense_large_input_t_layer2_t_config2_if_and_nl
      = IndexLoop_stage_0 & (~ IndexLoop_IndexLoop_nor_tmp);
  assign nnet_dense_large_input_t_layer2_t_config2_if_nnet_dense_large_input_t_layer2_t_config2_if_and_1_nl
      = IndexLoop_stage_0 & (~ (z_out_12[11]));
  assign and_830_nl = z_out_1_3 & IndexLoop_stage_0;
  assign IndexLoop_or_1_nl = and_dcpl_55 | (and_dcpl_100 & and_dcpl_517);
  assign IndexLoop_mux1h_9_nl = MUX1HOT_s_1_3_2((nnet_dense_large_input_t_layer2_t_config2_if_nnet_dense_large_input_t_layer2_t_config2_if_and_nl),
      (nnet_dense_large_input_t_layer2_t_config2_if_nnet_dense_large_input_t_layer2_t_config2_if_and_1_nl),
      (and_830_nl), {and_dcpl_65 , and_dcpl_60 , (IndexLoop_or_1_nl)});
  assign or_1413_nl = (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[4]) | (~
      (fsm_output[6])) | (fsm_output[7]);
  assign or_1414_nl = (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]);
  assign or_461_nl = (fsm_output[6]) | (fsm_output[3]) | (fsm_output[4]) | (~ (fsm_output[7]));
  assign mux_881_nl = MUX_s_1_2_2((or_1414_nl), (or_461_nl), fsm_output[2]);
  assign mux_882_nl = MUX_s_1_2_2((or_1413_nl), (mux_881_nl), fsm_output[1]);
  assign or_1416_nl = (fsm_output[1]) | (~ (fsm_output[2])) | (~ (fsm_output[3]))
      | (~ (fsm_output[4])) | (fsm_output[6]) | (~ (fsm_output[7]));
  assign mux_883_nl = MUX_s_1_2_2((mux_882_nl), (or_1416_nl), fsm_output[0]);
  assign mux_687_nl = MUX_s_1_2_2(or_tmp_91, or_864_cse, fsm_output[2]);
  assign mux_688_nl = MUX_s_1_2_2(or_381_cse, (mux_687_nl), fsm_output[1]);
  assign nl_IndexLoop_if_acc_nl = nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc14_sva_1
      + 6'b000001;
  assign IndexLoop_if_acc_nl = nl_IndexLoop_if_acc_nl[5:0];
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_and_14_nl
      = ((z_out_3!=6'b000000) | (z_out_13[3:0]!=4'b0000)) & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_mux_nl
      = MUX_v_6_2_2((IndexLoop_if_acc_nl), nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_5_0_pc14_sva_1,
      nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_outstep_and_14_nl);
  assign nor_217_nl = ~((~ (fsm_output[1])) | (fsm_output[2]) | (fsm_output[3]) |
      (fsm_output[4]) | (fsm_output[7]));
  assign mux_10_nl = MUX_s_1_2_2((~ or_tmp_2), and_2631_cse, fsm_output[3]);
  assign nor_353_nl = ~((fsm_output[1]) | (~((fsm_output[2]) & (mux_10_nl))));
  assign mux_890_nl = MUX_s_1_2_2((nor_217_nl), (nor_353_nl), fsm_output[0]);
  assign nand_148_nl = ~((mux_890_nl) & and_dcpl);
  assign or_1553_nl = (InitAccumLoop_1_iacc_6_0_sva_5_0[5]) | (fsm_output[2]) | (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]!=5'b00000)
      | (~ (fsm_output[1]));
  assign nand_158_nl = ~(IndexLoop_stage_0_2 & (~(and_2658_cse | (fsm_output[2])
      | (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]!=5'b00000) | (~ (fsm_output[1])))));
  assign mux_1054_nl = MUX_s_1_2_2((or_1553_nl), (nand_158_nl), fsm_output[0]);
  assign nand_213_nl = ~((fsm_output[0]) & IndexLoop_stage_0_2 & (fsm_output[2:1]==2'b10));
  assign mux_1055_nl = MUX_s_1_2_2((mux_1054_nl), (nand_213_nl), fsm_output[6]);
  assign or_1547_nl = (InitAccumLoop_2_iacc_3_0_sva!=4'b0000) | (~ and_817_cse);
  assign nand_157_nl = ~(IndexLoop_stage_0_2 & (~(and_2658_cse | (ReuseLoop_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_outidx_const_assign_1_ReuseLoop_2_asn_tmp_3_2_0_psp_sva_1!=3'b000)
      | (~ and_817_cse))));
  assign mux_1053_nl = MUX_s_1_2_2((or_1547_nl), (nand_157_nl), fsm_output[0]);
  assign or_1548_nl = (fsm_output[6]) | (mux_1053_nl);
  assign mux_1056_nl = MUX_s_1_2_2((mux_1055_nl), (or_1548_nl), fsm_output[7]);
  assign nor_663_nl = ~((fsm_output[4]) | (mux_1056_nl));
  assign nor_666_nl = ~((~ (fsm_output[7])) | (fsm_output[6]) | (fsm_output[2]) |
      (fsm_output[1]));
  assign mux_1051_nl = MUX_s_1_2_2(nor_668_cse, and_817_cse, fsm_output[0]);
  assign nor_667_nl = ~((fsm_output[7:6]!=2'b10) | (mux_1051_nl));
  assign mux_1052_nl = MUX_s_1_2_2((nor_666_nl), (nor_667_nl), fsm_output[4]);
  assign mux_1057_nl = MUX_s_1_2_2((nor_663_nl), (mux_1052_nl), fsm_output[3]);
  assign nor_669_nl = ~((InitAccumLoop_1_iacc_6_0_sva_5_0[5]) | (fsm_output[4]) |
      (fsm_output[2]) | (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]!=5'b00000) | (~ (fsm_output[1])));
  assign and_2660_nl = IndexLoop_stage_0_2 & (~(and_2658_cse | (fsm_output[4]) |
      (fsm_output[2]) | (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]!=5'b00000) | (~ (fsm_output[1]))));
  assign mux_1061_nl = MUX_s_1_2_2((nor_669_nl), (and_2660_nl), fsm_output[0]);
  assign nor_671_nl = ~((~ (fsm_output[0])) | (~ IndexLoop_stage_0_2) | (fsm_output[4])
      | (~ (fsm_output[2])) | (fsm_output[1]));
  assign mux_1062_nl = MUX_s_1_2_2((mux_1061_nl), (nor_671_nl), fsm_output[6]);
  assign or_1561_nl = (InitAccumLoop_2_iacc_3_0_sva!=4'b0000) | (fsm_output[4]) |
      nand_52_cse;
  assign nand_160_nl = ~(IndexLoop_stage_0_2 & (~(and_2658_cse | (ReuseLoop_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_outidx_const_assign_1_ReuseLoop_2_asn_tmp_3_2_0_psp_sva_1!=3'b000)
      | (fsm_output[4]) | nand_52_cse)));
  assign mux_1060_nl = MUX_s_1_2_2((or_1561_nl), (nand_160_nl), fsm_output[0]);
  assign nor_672_nl = ~((fsm_output[6]) | (mux_1060_nl));
  assign mux_1063_nl = MUX_s_1_2_2((mux_1062_nl), (nor_672_nl), fsm_output[7]);
  assign mux_1058_nl = MUX_s_1_2_2(or_10_cse, (~ or_10_cse), fsm_output[4]);
  assign nand_159_nl = ~((fsm_output[4]) & nand_52_cse);
  assign mux_1059_nl = MUX_s_1_2_2((mux_1058_nl), (nand_159_nl), fsm_output[0]);
  assign nor_674_nl = ~((fsm_output[7:6]!=2'b10) | (mux_1059_nl));
  assign mux_1064_nl = MUX_s_1_2_2((mux_1063_nl), (nor_674_nl), fsm_output[3]);
  assign nor_675_nl = ~((fsm_output[2]) | (InitAccumLoop_1_iacc_6_0_sva_5_0!=6'b000000)
      | (~ (fsm_output[1])) | (fsm_output[3]) | (fsm_output[6]));
  assign nor_676_nl = ~((InitAccumLoop_1_iacc_6_0_sva_5_0[4:0]!=5'b00000) | (~ (fsm_output[1]))
      | (fsm_output[3]) | (fsm_output[6]));
  assign nor_677_nl = ~((fsm_output[1]) | (fsm_output[3]) | (~ (fsm_output[6])));
  assign mux_1067_nl = MUX_s_1_2_2((nor_676_nl), (nor_677_nl), fsm_output[2]);
  assign nor_678_nl = ~((~ (fsm_output[2])) | (fsm_output[1]) | (fsm_output[3]) |
      (~ (fsm_output[6])));
  assign mux_1068_nl = MUX_s_1_2_2((mux_1067_nl), (nor_678_nl), and_2658_cse);
  assign and_2663_nl = IndexLoop_stage_0_2 & (mux_1068_nl);
  assign mux_1069_nl = MUX_s_1_2_2((nor_675_nl), (and_2663_nl), fsm_output[0]);
  assign nor_679_nl = ~((fsm_output[1]) | (~ (fsm_output[3])) | (fsm_output[6]));
  assign nor_680_nl = ~((InitAccumLoop_2_iacc_3_0_sva!=4'b0000) | (~ (fsm_output[1]))
      | (fsm_output[3]) | (fsm_output[6]));
  assign mux_1065_nl = MUX_s_1_2_2((nor_679_nl), (nor_680_nl), fsm_output[2]);
  assign and_2665_nl = IndexLoop_stage_0_2 & (~(and_2658_cse | (~ (fsm_output[2]))
      | (ReuseLoop_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer5_t_layer6_t_config6_outidx_const_assign_1_ReuseLoop_2_asn_tmp_3_2_0_psp_sva_1!=3'b000)
      | (~ (fsm_output[1])) | (fsm_output[3]) | (fsm_output[6])));
  assign mux_1066_nl = MUX_s_1_2_2((mux_1065_nl), (and_2665_nl), fsm_output[0]);
  assign mux_1070_nl = MUX_s_1_2_2((mux_1069_nl), (mux_1066_nl), fsm_output[7]);
  assign nor_682_nl = ~((~ (fsm_output[7])) | (~ (fsm_output[0])) | (fsm_output[2])
      | (fsm_output[1]) | (~ (fsm_output[3])) | (fsm_output[6]));
  assign mux_1071_nl = MUX_s_1_2_2((mux_1070_nl), (nor_682_nl), fsm_output[4]);
  assign and_591_nl = and_dcpl_588 & and_dcpl_587;
  assign and_593_nl = and_dcpl_590 & and_dcpl_587;
  assign mux_934_nl = MUX_s_1_2_2(mux_tmp_933, mux_tmp_500, fsm_output[0]);
  assign and_587_nl = and_dcpl_64 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_482_m1c;
  assign and_588_nl = and_dcpl_59 & and_dcpl_584;
  assign mux_522_nl = MUX_s_1_2_2(mux_tmp_521, mux_tmp_519, fsm_output[1]);
  assign mux_523_nl = MUX_s_1_2_2((mux_522_nl), mux_tmp_520, fsm_output[0]);
  assign nor_659_nl = ~((fsm_output[2:0]!=3'b011) | (~ IndexLoop_stage_0_2) | (fsm_output[3]));
  assign nor_660_nl = ~((fsm_output[2:0]!=3'b101) | IndexLoop_stage_0 | (~ IndexLoop_stage_0_2)
      | (fsm_output[3]));
  assign mux_1072_nl = MUX_s_1_2_2((nor_659_nl), (nor_660_nl), fsm_output[6]);
  assign nor_661_nl = ~((fsm_output[6]) | and_2657_cse | (~ (fsm_output[3])));
  assign mux_1073_nl = MUX_s_1_2_2((mux_1072_nl), (nor_661_nl), fsm_output[7]);
  assign mux_1074_nl = MUX_s_1_2_2((mux_1073_nl), nor_662_cse, fsm_output[4]);
  assign nor_655_nl = ~((~ IndexLoop_stage_0_2) | (fsm_output[2]) | (~ (fsm_output[1]))
      | (fsm_output[7]) | (~ (fsm_output[0])));
  assign nor_656_nl = ~((fsm_output[2]) | (fsm_output[1]) | (~ (fsm_output[7])) |
      (fsm_output[0]));
  assign mux_1075_nl = MUX_s_1_2_2((nor_655_nl), (nor_656_nl), fsm_output[3]);
  assign nor_657_nl = ~((fsm_output[3]) | (~ IndexLoop_stage_0_2) | (fsm_output[2:1]!=2'b10)
      | IndexLoop_stage_0 | (fsm_output[7]) | (~ (fsm_output[0])));
  assign mux_1076_nl = MUX_s_1_2_2((mux_1075_nl), (nor_657_nl), fsm_output[6]);
  assign mux_1077_nl = MUX_s_1_2_2((mux_1076_nl), nor_662_cse, fsm_output[4]);
  assign and_638_nl = and_dcpl_624 & and_dcpl_57;
  assign and_639_nl = and_dcpl_626 & and_dcpl_57;
  assign and_662_nl = and_dcpl_659 & and_dcpl_587;
  assign and_664_nl = and_dcpl_661 & and_dcpl_587;
  assign mux_950_nl = MUX_s_1_2_2(mux_tmp_738, mux_tmp_774, fsm_output[0]);
  assign and_685_nl = and_dcpl_659 & and_dcpl_573;
  assign and_686_nl = and_dcpl_661 & and_dcpl_573;
  assign and_705_nl = and_dcpl_59 & and_dcpl_62;
  assign and_709_nl = and_dcpl_54 & and_dcpl_62;
  assign and_702_nl = and_dcpl_59 & and_dcpl_154;
  assign and_704_nl = and_dcpl_54 & and_dcpl_154;
  assign mux_959_nl = MUX_s_1_2_2(mux_425_cse, mux_tmp_419, fsm_output[0]);
  assign and_595_nl = and_dcpl_588 & and_dcpl_592;
  assign and_596_nl = and_dcpl_590 & and_dcpl_592;
  assign and_699_nl = and_dcpl_59 & and_dcpl_592;
  assign and_701_nl = and_dcpl_54 & and_dcpl_592;
  assign and_696_nl = and_dcpl_59 & and_dcpl_587;
  assign and_698_nl = and_dcpl_54 & and_dcpl_587;
  assign mux_417_nl = MUX_s_1_2_2(mux_661_cse, or_864_cse, and_817_cse);
  assign mux_958_nl = MUX_s_1_2_2(mux_tmp_419, (mux_417_nl), fsm_output[0]);
  assign and_693_nl = and_dcpl_659 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_472_m1c;
  assign and_695_nl = and_dcpl_661 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_472_m1c;
  assign and_691_nl = and_dcpl_659 & and_dcpl_517;
  assign and_692_nl = and_dcpl_661 & and_dcpl_517;
  assign mux_957_nl = MUX_s_1_2_2(mux_tmp_587, mux_tmp_594, fsm_output[0]);
  assign mux_171_nl = MUX_s_1_2_2(mux_661_cse, or_864_cse, fsm_output[1]);
  assign or_870_nl = (fsm_output[1]) | (fsm_output[6]) | (~ (fsm_output[7]));
  assign mux_603_nl = MUX_s_1_2_2((mux_171_nl), (or_870_nl), fsm_output[0]);
  assign mux_604_nl = MUX_s_1_2_2(mux_661_cse, (mux_603_nl), fsm_output[2]);
  assign or_1001_nl = nor_668_cse | (fsm_output[7]);
  assign mux_605_nl = MUX_s_1_2_2((mux_604_nl), (or_1001_nl), fsm_output[4]);
  assign or_649_nl = (~ (fsm_output[4])) | (fsm_output[7]);
  assign mux_606_nl = MUX_s_1_2_2((mux_605_nl), (or_649_nl), fsm_output[3]);
  assign mux_607_nl = MUX_s_1_2_2((mux_606_nl), (fsm_output[7]), fsm_output[5]);
  assign or_1598_nl = and_2654_cse | (fsm_output[4:3]!=2'b10);
  assign mux_1080_nl = MUX_s_1_2_2((or_1598_nl), or_tmp_922, fsm_output[0]);
  assign nand_164_nl = ~((fsm_output[1]) & (~ (mux_1080_nl)));
  assign or_1596_nl = (fsm_output[1]) | (~ (fsm_output[0])) | (~ (fsm_output[6]))
      | (fsm_output[3]) | IndexLoop_stage_0 | (~ IndexLoop_stage_0_2) | (fsm_output[4]);
  assign mux_1081_nl = MUX_s_1_2_2((nand_164_nl), (or_1596_nl), fsm_output[2]);
  assign or_1595_nl = (~ (fsm_output[1])) | (fsm_output[6]) | not_tmp_1409;
  assign or_1593_nl = (fsm_output[6]) | not_tmp_1409;
  assign mux_1078_nl = MUX_s_1_2_2((or_1593_nl), or_tmp_922, and_810_cse_1);
  assign mux_1079_nl = MUX_s_1_2_2((or_1595_nl), (mux_1078_nl), fsm_output[2]);
  assign mux_1082_nl = MUX_s_1_2_2((mux_1081_nl), (mux_1079_nl), fsm_output[7]);
  assign nor_650_nl = ~((fsm_output[2:0]!=3'b101));
  assign mux_1084_nl = MUX_s_1_2_2(nor_649_cse, (nor_650_nl), fsm_output[6]);
  assign nor_651_nl = ~((fsm_output[6]) | nand_210_cse);
  assign mux_1085_nl = MUX_s_1_2_2((mux_1084_nl), (nor_651_nl), fsm_output[7]);
  assign and_2656_nl = (~(IndexLoop_stage_0 | (~ IndexLoop_stage_0_2))) & (mux_1085_nl);
  assign nor_652_nl = ~((fsm_output[7]) | (fsm_output[2]) | (~ (fsm_output[1])) |
      (fsm_output[0]));
  assign nor_653_nl = ~((fsm_output[7]) | (fsm_output[6]) | (fsm_output[2]) | (~
      (fsm_output[1])) | (fsm_output[0]));
  assign mux_1083_nl = MUX_s_1_2_2((nor_652_nl), (nor_653_nl), z_out_23_22_8[10]);
  assign mux_1086_nl = MUX_s_1_2_2((and_2656_nl), (mux_1083_nl), fsm_output[4]);
  assign mux_1087_nl = MUX_s_1_2_2((mux_1086_nl), nor_654_cse, fsm_output[3]);
  assign ReuseLoop_ReuseLoop_and_nl = (z_out_2[9:0]) & (signext_10_1(z_out_11[7]))
      & ({{9{and_dcpl_65}}, and_dcpl_65});
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_470_nl =
      and_dcpl_155 | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_566_rgt;
  assign nor_945_nl = ~((fsm_output[7:6]!=2'b01) | IndexLoop_stage_0 | (~ IndexLoop_stage_0_2)
      | (fsm_output[4]) | not_tmp_1420);
  assign nor_946_nl = ~((or_1876_cse & (fsm_output[0])) | (fsm_output[2]));
  assign nor_947_nl = ~((z_out_23_22_8[10]) | (~ (fsm_output[4])) | (fsm_output[0])
      | (fsm_output[2]));
  assign mux_1088_nl = MUX_s_1_2_2((nor_946_nl), (nor_947_nl), fsm_output[6]);
  assign nor_948_nl = ~((fsm_output[6]) | IndexLoop_stage_0 | (~ IndexLoop_stage_0_2)
      | (fsm_output[4]) | not_tmp_1420);
  assign mux_1089_nl = MUX_s_1_2_2((mux_1088_nl), (nor_948_nl), fsm_output[7]);
  assign mux_1090_nl = MUX_s_1_2_2((nor_945_nl), (mux_1089_nl), fsm_output[1]);
  assign mux_1091_nl = MUX_s_1_2_2((mux_1090_nl), nor_654_cse, fsm_output[3]);
  assign and_689_nl = and_dcpl_659 & and_dcpl_579;
  assign and_690_nl = and_dcpl_661 & and_dcpl_579;
  assign mux_435_nl = MUX_s_1_2_2(mux_tmp_81, or_tmp_48, or_647_cse_1);
  assign mux_621_nl = MUX_s_1_2_2(mux_tmp_620, (mux_435_nl), fsm_output[1]);
  assign mux_623_nl = MUX_s_1_2_2(mux_tmp_622, (mux_621_nl), fsm_output[0]);
  assign or_1623_nl = (fsm_output[7]) | (fsm_output[2]) | (~ and_810_cse_1);
  assign mux_1097_nl = MUX_s_1_2_2(nand_tmp_52, (or_1623_nl), fsm_output[4]);
  assign mux_1096_nl = MUX_s_1_2_2(nand_tmp_52, or_tmp_948, fsm_output[4]);
  assign mux_1098_nl = MUX_s_1_2_2((mux_1097_nl), (mux_1096_nl), z_out_23_22_8[10]);
  assign mux_1092_nl = MUX_s_1_2_2((~ and_810_cse_1), and_810_cse_1, fsm_output[2]);
  assign or_1616_nl = (~ (fsm_output[4])) | (~ (fsm_output[7])) | (fsm_output[6])
      | (mux_1092_nl);
  assign mux_1099_nl = MUX_s_1_2_2((mux_1098_nl), (or_1616_nl), fsm_output[3]);
  assign or_1632_nl = (fsm_output[7]) | (fsm_output[2]) | (~ (fsm_output[1]));
  assign mux_1104_nl = MUX_s_1_2_2(nand_tmp_53, (or_1632_nl), fsm_output[4]);
  assign mux_1103_nl = MUX_s_1_2_2(nand_tmp_53, or_tmp_957, fsm_output[4]);
  assign mux_1105_nl = MUX_s_1_2_2((mux_1104_nl), (mux_1103_nl), z_out_23_22_8[10]);
  assign or_1625_nl = (~ (fsm_output[4])) | (~ (fsm_output[7])) | (fsm_output[6])
      | (fsm_output[2]) | (~ (fsm_output[1]));
  assign mux_1106_nl = MUX_s_1_2_2((mux_1105_nl), (or_1625_nl), fsm_output[3]);
  assign and_687_nl = and_dcpl_659 & and_dcpl_576;
  assign and_688_nl = and_dcpl_661 & and_dcpl_576;
  assign mux_956_nl = MUX_s_1_2_2(mux_tmp_594, mux_tmp_555, fsm_output[0]);
  assign mux_636_nl = MUX_s_1_2_2(mux_tmp_622, mux_tmp_635, fsm_output[0]);
  assign nor_641_nl = ~((fsm_output[0]) | (fsm_output[3]) | (~ (fsm_output[2])));
  assign mux_1110_nl = MUX_s_1_2_2((nor_641_nl), and_2650_cse, fsm_output[7]);
  assign and_2651_nl = (fsm_output[4]) & (mux_1110_nl);
  assign nor_643_nl = ~((z_out_23_22_8[10]) | (fsm_output[7]) | (fsm_output[0]) |
      (fsm_output[3]) | (~ (fsm_output[2])));
  assign mux_1109_nl = MUX_s_1_2_2(nor_642_cse, (nor_643_nl), fsm_output[4]);
  assign mux_1111_nl = MUX_s_1_2_2((and_2651_nl), (mux_1109_nl), fsm_output[6]);
  assign or_1636_nl = (~ (fsm_output[0])) | (~ IndexLoop_stage_0_2) | IndexLoop_stage_0
      | (fsm_output[3:2]!=2'b01);
  assign mux_1107_nl = MUX_s_1_2_2(or_1637_cse, (or_1636_nl), fsm_output[7]);
  assign or_1634_nl = (~ (fsm_output[7])) | (fsm_output[0]) | (~ and_2650_cse);
  assign mux_1108_nl = MUX_s_1_2_2((mux_1107_nl), (or_1634_nl), fsm_output[4]);
  assign nor_644_nl = ~((fsm_output[6]) | (mux_1108_nl));
  assign mux_1112_nl = MUX_s_1_2_2((mux_1111_nl), (nor_644_nl), fsm_output[1]);
  assign or_1656_nl = (~ (fsm_output[4])) | (fsm_output[0]) | (~ (fsm_output[2]));
  assign nand_214_nl = ~((fsm_output[0]) & IndexLoop_stage_0_2 & (~ IndexLoop_stage_0)
      & (fsm_output[2]));
  assign or_1652_nl = (fsm_output[0]) | (~ (fsm_output[2]));
  assign mux_1114_nl = MUX_s_1_2_2((nand_214_nl), (or_1652_nl), fsm_output[4]);
  assign or_1651_nl = (fsm_output[4]) | (~ (fsm_output[0])) | (~ IndexLoop_stage_0_2)
      | IndexLoop_stage_0 | (~ (fsm_output[2]));
  assign mux_1115_nl = MUX_s_1_2_2((mux_1114_nl), (or_1651_nl), z_out_23_22_8[10]);
  assign mux_1116_nl = MUX_s_1_2_2((or_1656_nl), (mux_1115_nl), fsm_output[6]);
  assign nor_645_nl = ~((fsm_output[7]) | (mux_1116_nl));
  assign mux_1113_nl = MUX_s_1_2_2(nor_646_cse, nor_647_cse, fsm_output[7]);
  assign mux_1117_nl = MUX_s_1_2_2((nor_645_nl), (mux_1113_nl), fsm_output[1]);
  assign nor_648_nl = ~((fsm_output[1]) | (~ (fsm_output[7])) | (fsm_output[6]) |
      (~ (fsm_output[4])) | (fsm_output[0]) | (~ (fsm_output[2])));
  assign mux_1118_nl = MUX_s_1_2_2((mux_1117_nl), (nor_648_nl), fsm_output[3]);
  assign and_683_nl = and_dcpl_659 & and_dcpl_570;
  assign and_684_nl = and_dcpl_661 & and_dcpl_570;
  assign mux_955_nl = MUX_s_1_2_2(mux_tmp_555, mux_tmp_642, fsm_output[0]);
  assign mux_647_nl = MUX_s_1_2_2(mux_tmp_646, mux_tmp_635, fsm_output[0]);
  assign nor_633_nl = ~((fsm_output[3]) | not_tmp_1420);
  assign and_2649_nl = (fsm_output[3]) & (fsm_output[2]) & (fsm_output[0]);
  assign mux_1122_nl = MUX_s_1_2_2((nor_633_nl), (and_2649_nl), fsm_output[7]);
  assign and_2648_nl = (fsm_output[4]) & (mux_1122_nl);
  assign nor_634_nl = ~((fsm_output[7]) | (~ IndexLoop_stage_0_2) | IndexLoop_stage_0
      | (fsm_output[3]) | not_tmp_1420);
  assign nor_635_nl = ~((z_out_23_22_8[10]) | (fsm_output[7]) | (fsm_output[3]) |
      not_tmp_1420);
  assign mux_1121_nl = MUX_s_1_2_2((nor_634_nl), (nor_635_nl), fsm_output[4]);
  assign mux_1123_nl = MUX_s_1_2_2((and_2648_nl), (mux_1121_nl), fsm_output[6]);
  assign or_1660_nl = (~ IndexLoop_stage_0_2) | IndexLoop_stage_0 | (fsm_output[3])
      | not_tmp_1420;
  assign mux_1119_nl = MUX_s_1_2_2(or_1637_cse, (or_1660_nl), fsm_output[7]);
  assign nand_204_nl = ~((fsm_output[7]) & (fsm_output[3]) & (fsm_output[2]) & (~
      (fsm_output[0])));
  assign mux_1120_nl = MUX_s_1_2_2((mux_1119_nl), (nand_204_nl), fsm_output[4]);
  assign nor_636_nl = ~((fsm_output[6]) | (mux_1120_nl));
  assign mux_1124_nl = MUX_s_1_2_2((mux_1123_nl), (nor_636_nl), fsm_output[1]);
  assign nor_637_nl = ~((fsm_output[7:6]!=2'b01) | (~ IndexLoop_stage_0_2) | IndexLoop_stage_0
      | (fsm_output[3:2]!=2'b01));
  assign nor_638_nl = ~((fsm_output[3:2]!=2'b01));
  assign mux_1126_nl = MUX_s_1_2_2((nor_638_nl), and_2650_cse, fsm_output[7]);
  assign nor_639_nl = ~((z_out_23_22_8[10]) | (fsm_output[7]) | (fsm_output[3]) |
      (~ (fsm_output[2])));
  assign mux_1127_nl = MUX_s_1_2_2((mux_1126_nl), (nor_639_nl), fsm_output[6]);
  assign mux_1128_nl = MUX_s_1_2_2((nor_637_nl), (mux_1127_nl), fsm_output[4]);
  assign or_1672_nl = (~ IndexLoop_stage_0_2) | (fsm_output[3:2]!=2'b00);
  assign or_1671_nl = (~ IndexLoop_stage_0_2) | IndexLoop_stage_0 | (fsm_output[3:2]!=2'b01);
  assign mux_1125_nl = MUX_s_1_2_2((or_1672_nl), (or_1671_nl), fsm_output[7]);
  assign nor_640_nl = ~((fsm_output[4]) | (fsm_output[6]) | (mux_1125_nl));
  assign mux_1129_nl = MUX_s_1_2_2((mux_1128_nl), (nor_640_nl), fsm_output[1]);
  assign and_681_nl = and_dcpl_659 & and_dcpl_567;
  assign and_682_nl = and_dcpl_661 & and_dcpl_567;
  assign mux_658_nl = MUX_s_1_2_2(mux_tmp_646, mux_tmp_657, fsm_output[0]);
  assign and_605_nl = and_dcpl_588 & and_dcpl_159;
  assign and_606_nl = and_dcpl_590 & and_dcpl_159;
  assign nor_954_nl = ~((fsm_output[7]) | (~ (fsm_output[6])) | (~ (fsm_output[2]))
      | IndexLoop_stage_0 | (~ IndexLoop_stage_0_2) | (fsm_output[4]) | (~ (fsm_output[0])));
  assign nor_955_nl = ~((~ IndexLoop_stage_0_2) | (fsm_output[4]) | (~ (fsm_output[0])));
  assign nor_956_nl = ~((~ (fsm_output[4])) | (fsm_output[0]));
  assign mux_1130_nl = MUX_s_1_2_2((nor_955_nl), (nor_956_nl), fsm_output[2]);
  assign nor_957_nl = ~((z_out_23_22_8[10]) | (~ (fsm_output[2])) | (~ (fsm_output[4]))
      | (fsm_output[0]));
  assign mux_1131_nl = MUX_s_1_2_2((mux_1130_nl), (nor_957_nl), fsm_output[6]);
  assign mux_1132_nl = MUX_s_1_2_2((mux_1131_nl), nor_647_cse, fsm_output[7]);
  assign mux_1133_nl = MUX_s_1_2_2((nor_954_nl), (mux_1132_nl), fsm_output[1]);
  assign and_679_nl = and_dcpl_659 & and_dcpl_519;
  assign and_680_nl = and_dcpl_661 & and_dcpl_519;
  assign mux_954_nl = MUX_s_1_2_2(mux_tmp_642, mux_tmp_680, fsm_output[0]);
  assign mux_671_nl = MUX_s_1_2_2(mux_tmp_670, mux_tmp_657, fsm_output[0]);
  assign and_607_nl = and_dcpl_588 & and_dcpl_51;
  assign and_608_nl = and_dcpl_590 & and_dcpl_51;
  assign or_1694_nl = (fsm_output[7]) | nand_52_cse;
  assign mux_1138_nl = MUX_s_1_2_2(nand_tmp_54, (or_1694_nl), fsm_output[4]);
  assign or_1688_nl = (fsm_output[7:6]!=2'b00) | nand_52_cse;
  assign mux_1137_nl = MUX_s_1_2_2(nand_tmp_54, (or_1688_nl), fsm_output[4]);
  assign mux_1139_nl = MUX_s_1_2_2((mux_1138_nl), (mux_1137_nl), z_out_23_22_8[10]);
  assign and_677_nl = and_dcpl_659 & and_dcpl_51;
  assign and_678_nl = and_dcpl_661 & and_dcpl_51;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_259_nl =
      (and_dcpl_334 & and_dcpl_261 & and_dcpl_65) | (and_dcpl_189 & (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_out_index_4_0_sva_1[4])
      & and_dcpl_227 & and_dcpl_60) | ((~ or_1084_tmp) & and_dcpl_55);
  assign MultLoop_and_181_nl = (~ or_dcpl_599) & and_397_m1c & and_dcpl_65;
  assign MultLoop_and_182_nl = or_dcpl_599 & and_397_m1c & and_dcpl_65;
  assign and_400_nl = or_dcpl_522 & IndexLoop_stage_0_2 & and_dcpl_60;
  assign and_675_nl = and_dcpl_659 & and_dcpl_159;
  assign and_676_nl = and_dcpl_661 & and_dcpl_159;
  assign mux_953_nl = MUX_s_1_2_2(mux_tmp_680, mux_tmp_691, fsm_output[0]);
  assign mux_698_nl = MUX_s_1_2_2(mux_tmp_521, mux_tmp_517, or_1875_cse);
  assign nor_623_nl = ~((~ (fsm_output[7])) | (fsm_output[4]) | (~ (fsm_output[3]))
      | (fsm_output[6]) | (fsm_output[2]));
  assign nor_624_nl = ~((fsm_output[3]) | (~ (fsm_output[6])) | IndexLoop_stage_0
      | (~ (fsm_output[2])));
  assign nor_625_nl = ~((fsm_output[3]) | (fsm_output[6]) | (fsm_output[2]));
  assign mux_1141_nl = MUX_s_1_2_2((nor_624_nl), (nor_625_nl), fsm_output[1]);
  assign and_2647_nl = IndexLoop_stage_0_2 & (mux_1141_nl);
  assign nor_626_nl = ~((fsm_output[3:1]!=3'b100));
  assign nor_627_nl = ~((fsm_output[1]) | (~ (fsm_output[3])) | (fsm_output[6]) |
      (fsm_output[2]));
  assign mux_1140_nl = MUX_s_1_2_2((nor_626_nl), (nor_627_nl), z_out_23_22_8[10]);
  assign mux_1142_nl = MUX_s_1_2_2((and_2647_nl), (mux_1140_nl), fsm_output[4]);
  assign nor_628_nl = ~((fsm_output[4]) | (fsm_output[1]) | (~ (fsm_output[3])) |
      (fsm_output[6]) | (fsm_output[2]));
  assign mux_1143_nl = MUX_s_1_2_2((mux_1142_nl), (nor_628_nl), fsm_output[7]);
  assign mux_1144_nl = MUX_s_1_2_2((nor_623_nl), (mux_1143_nl), fsm_output[0]);
  assign nor_619_nl = ~((fsm_output[3:1]!=3'b001));
  assign nor_620_nl = ~((fsm_output[3:2]!=2'b01) | IndexLoop_stage_0 | (fsm_output[1]));
  assign mux_1145_nl = MUX_s_1_2_2((nor_619_nl), (nor_620_nl), fsm_output[6]);
  assign and_2645_nl = IndexLoop_stage_0_2 & (mux_1145_nl);
  assign nor_621_nl = ~(and_2654_cse | (fsm_output[3:1]!=3'b100));
  assign mux_1146_nl = MUX_s_1_2_2((and_2645_nl), (nor_621_nl), fsm_output[4]);
  assign and_2644_nl = (fsm_output[0]) & (mux_1146_nl);
  assign mux_1147_nl = MUX_s_1_2_2((and_2644_nl), nor_622_cse, fsm_output[7]);
  assign and_673_nl = and_dcpl_659 & and_dcpl_57;
  assign and_674_nl = and_dcpl_661 & and_dcpl_57;
  assign mux_708_nl = MUX_s_1_2_2(mux_tmp_707, mux_tmp_520, fsm_output[0]);
  assign nor_615_nl = ~((fsm_output[3]) | (~ (fsm_output[0])) | (~ IndexLoop_stage_0_2)
      | (fsm_output[4]) | (~ (fsm_output[6])) | IndexLoop_stage_0 | (~ (fsm_output[2])));
  assign nor_617_nl = ~((fsm_output[0]) | (~ (fsm_output[4])) | (fsm_output[2]));
  assign mux_1148_nl = MUX_s_1_2_2(nor_646_cse, (nor_617_nl), fsm_output[3]);
  assign mux_1149_nl = MUX_s_1_2_2((nor_615_nl), (mux_1148_nl), fsm_output[1]);
  assign nor_618_nl = ~((~ (fsm_output[3])) | (fsm_output[4]) | (fsm_output[6]) |
      (fsm_output[2]));
  assign mux_1150_nl = MUX_s_1_2_2((mux_1149_nl), (nor_618_nl), fsm_output[7]);
  assign nor_611_nl = ~((fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[3]))
      | (fsm_output[0]));
  assign mux_1151_nl = MUX_s_1_2_2((nor_611_nl), nor_642_cse, fsm_output[6]);
  assign nor_613_nl = ~((fsm_output[6]) | (fsm_output[2]) | (fsm_output[7]) | (~
      IndexLoop_stage_0_2) | (fsm_output[3]) | (~ (fsm_output[0])));
  assign mux_1152_nl = MUX_s_1_2_2((mux_1151_nl), (nor_613_nl), fsm_output[1]);
  assign nor_614_nl = ~((~ (fsm_output[1])) | (fsm_output[2]) | (fsm_output[7]) |
      (~ (fsm_output[3])) | (fsm_output[0]));
  assign mux_1153_nl = MUX_s_1_2_2((mux_1152_nl), (nor_614_nl), fsm_output[4]);
  assign and_671_nl = and_dcpl_659 & and_dcpl_157;
  assign and_672_nl = and_dcpl_661 & and_dcpl_157;
  assign mux_952_nl = MUX_s_1_2_2(mux_tmp_691, mux_tmp_724, fsm_output[0]);
  assign mux_717_nl = MUX_s_1_2_2(mux_tmp_521, mux_tmp_519, or_1875_cse);
  assign and_2643_nl = (fsm_output[7]) & (fsm_output[3]);
  assign mux_1155_nl = MUX_s_1_2_2((and_2643_nl), nor_642_cse, fsm_output[6]);
  assign nor_609_nl = ~((~ IndexLoop_stage_0_2) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign mux_1154_nl = MUX_s_1_2_2((nor_609_nl), (fsm_output[3]), fsm_output[7]);
  assign nor_608_nl = ~((fsm_output[6]) | (fsm_output[2]) | (~ (mux_1154_nl)));
  assign mux_1156_nl = MUX_s_1_2_2((mux_1155_nl), (nor_608_nl), fsm_output[1]);
  assign mux_1157_nl = MUX_s_1_2_2((mux_1156_nl), nor_610_cse, fsm_output[4]);
  assign or_1729_nl = (~ (fsm_output[7])) | (~ (fsm_output[3])) | (fsm_output[0]);
  assign or_1728_nl = (~ IndexLoop_stage_0_2) | (fsm_output[7]) | (fsm_output[3])
      | (~ (fsm_output[0]));
  assign mux_1158_nl = MUX_s_1_2_2((or_1729_nl), (or_1728_nl), fsm_output[1]);
  assign nor_604_nl = ~((fsm_output[6]) | (mux_1158_nl));
  assign nor_605_nl = ~(IndexLoop_stage_0 | (~ (fsm_output[6])) | (fsm_output[1])
      | (~ IndexLoop_stage_0_2) | (fsm_output[7]) | (fsm_output[3]) | (~ (fsm_output[0])));
  assign mux_1159_nl = MUX_s_1_2_2((nor_604_nl), (nor_605_nl), fsm_output[2]);
  assign mux_1160_nl = MUX_s_1_2_2((mux_1159_nl), nor_610_cse, fsm_output[4]);
  assign and_669_nl = and_dcpl_659 & and_dcpl_62;
  assign and_670_nl = and_dcpl_661 & and_dcpl_62;
  assign mux_729_nl = MUX_s_1_2_2(mux_tmp_184, mux_tmp_513, and_2657_cse);
  assign nor_603_nl = ~((~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[4]) |
      and_2642_cse);
  assign mux_1163_nl = MUX_s_1_2_2(mux_1162_cse, (nor_603_nl), fsm_output[7]);
  assign mux_1166_nl = MUX_s_1_2_2(mux_1162_cse, nor_622_cse, fsm_output[7]);
  assign and_667_nl = and_dcpl_659 & and_dcpl_154;
  assign and_668_nl = and_dcpl_661 & and_dcpl_154;
  assign mux_951_nl = MUX_s_1_2_2(mux_tmp_724, mux_tmp_738, fsm_output[0]);
  assign mux_744_nl = MUX_s_1_2_2(mux_tmp_184, mux_tmp_513, and_817_cse);
  assign mux_743_nl = MUX_s_1_2_2(mux_tmp_742, mux_tmp_519, fsm_output[1]);
  assign mux_745_nl = MUX_s_1_2_2((mux_744_nl), (mux_743_nl), fsm_output[0]);
  assign nor_594_nl = ~((fsm_output[3:0]!=4'b0011));
  assign nor_595_nl = ~(IndexLoop_stage_0 | (fsm_output[3:0]!=4'b0101));
  assign mux_1167_nl = MUX_s_1_2_2((nor_594_nl), (nor_595_nl), fsm_output[6]);
  assign and_2637_nl = IndexLoop_stage_0_2 & (mux_1167_nl);
  assign nor_596_nl = ~((fsm_output[6]) | (~ (fsm_output[3])));
  assign mux_1168_nl = MUX_s_1_2_2((and_2637_nl), (nor_596_nl), fsm_output[7]);
  assign nor_597_nl = ~((fsm_output[7]) | (fsm_output[0]) | (~((fsm_output[3:1]==3'b111))));
  assign mux_1169_nl = MUX_s_1_2_2((mux_1168_nl), (nor_597_nl), fsm_output[4]);
  assign nor_589_nl = ~((fsm_output[2]) | (fsm_output[4]) | (~ (fsm_output[7])) |
      (~ (fsm_output[3])) | (fsm_output[0]));
  assign nor_590_nl = ~((~ (fsm_output[2])) | IndexLoop_stage_0 | (fsm_output[4])
      | (fsm_output[7]) | (~ IndexLoop_stage_0_2) | (fsm_output[3]) | (~ (fsm_output[0])));
  assign mux_1172_nl = MUX_s_1_2_2((nor_589_nl), (nor_590_nl), fsm_output[6]);
  assign nor_591_nl = ~((fsm_output[4]) | (fsm_output[7]) | (~ IndexLoop_stage_0_2)
      | (fsm_output[3]) | (~ (fsm_output[0])));
  assign nor_592_nl = ~((~ (fsm_output[4])) | (fsm_output[7]) | (~ (fsm_output[3]))
      | (fsm_output[0]));
  assign mux_1170_nl = MUX_s_1_2_2((nor_591_nl), (nor_592_nl), fsm_output[2]);
  assign nor_593_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[4])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[0]));
  assign mux_1171_nl = MUX_s_1_2_2((mux_1170_nl), (nor_593_nl), fsm_output[6]);
  assign mux_1173_nl = MUX_s_1_2_2((mux_1172_nl), (mux_1171_nl), fsm_output[1]);
  assign and_665_nl = and_dcpl_659 & and_dcpl_592;
  assign and_666_nl = and_dcpl_661 & and_dcpl_592;
  assign MultLoop_1_1_MultLoop_1_mux_nl = MUX_v_2_64_2(layer3_out_0_16_0_lpi_1_dfm_16_15,
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_16_0_lpi_1_dfm_16_12[4:3]),
      reg_nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_16_0_lpi_1_dfm_ftd,
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_16_0_lpi_1_dfm[16:15]),
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_16_0_lpi_1_dfm[16:15]),
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_16_0_lpi_1_dfm[16:15]),
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_16_0_lpi_1_dfm[16:15]),
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_16_0_lpi_1_dfm[16:15]),
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_16_0_lpi_1_dfm[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_63_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_2_reg[4:3]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_2_reg[4:3]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_2_reg[4:3]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_2_reg[4:3]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd_1[16:15]),
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_16_0_lpi_1_dfm[16:15]),
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_16_15,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_16_15,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_16_15,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_16_15,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_16_15,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_16_15,
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_16_0_lpi_1_dfm[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_1_ftd_1[16:15]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_1_ftd_1[16:15]),
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_16_0_lpi_1_dfm[16:15]),
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_16_0_lpi_1_dfm[16:15]),
      InitAccumLoop_1_iacc_6_0_sva_5_0);
  assign or_1771_nl = (~ (fsm_output[1])) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]);
  assign or_1770_nl = (~((~ (fsm_output[1])) | (fsm_output[4]))) | (fsm_output[7:6]!=2'b10);
  assign mux_1179_nl = MUX_s_1_2_2((or_1771_nl), (or_1770_nl), fsm_output[3]);
  assign or_1767_nl = (~ or_tmp_940) | (~ (fsm_output[1])) | (fsm_output[4]) | (fsm_output[6])
      | (fsm_output[7]);
  assign mux_1178_nl = MUX_s_1_2_2((or_1767_nl), or_tmp_1095, fsm_output[3]);
  assign mux_1180_nl = MUX_s_1_2_2((mux_1179_nl), (mux_1178_nl), fsm_output[0]);
  assign or_1763_nl = (~((fsm_output[1]) | (fsm_output[4]))) | (fsm_output[7:6]!=2'b10);
  assign or_1758_nl = (fsm_output[1]) | (fsm_output[4]);
  assign mux_1174_nl = MUX_s_1_2_2(or_865_cse_1, or_864_cse, or_1758_nl);
  assign mux_1175_nl = MUX_s_1_2_2((or_1763_nl), (mux_1174_nl), or_tmp_940);
  assign or_1756_nl = (fsm_output[1]) | (~ (fsm_output[4])) | (fsm_output[6]) | (~
      (fsm_output[7]));
  assign mux_1176_nl = MUX_s_1_2_2((mux_1175_nl), (or_1756_nl), fsm_output[3]);
  assign mux_1177_nl = MUX_s_1_2_2(or_tmp_1095, (mux_1176_nl), fsm_output[0]);
  assign mux_1181_nl = MUX_s_1_2_2((mux_1180_nl), (mux_1177_nl), fsm_output[2]);
  assign nor_583_nl = ~((~ (fsm_output[1])) | (fsm_output[6]) | (fsm_output[7]));
  assign and_2635_nl = (fsm_output[1]) & (~((~ or_tmp_940) | (fsm_output[7:6]!=2'b00)));
  assign mux_1183_nl = MUX_s_1_2_2((nor_583_nl), (and_2635_nl), fsm_output[0]);
  assign nor_585_nl = ~((~ or_tmp_940) | (fsm_output[7:6]!=2'b01));
  assign mux_1182_nl = MUX_s_1_2_2((nor_585_nl), nor_586_cse, fsm_output[1]);
  assign and_2636_nl = (fsm_output[0]) & (mux_1182_nl);
  assign mux_1184_nl = MUX_s_1_2_2((mux_1183_nl), (and_2636_nl), fsm_output[2]);
  assign nor_587_nl = ~((~ (fsm_output[2])) | (fsm_output[0]) | (fsm_output[1]) |
      (fsm_output[6]) | (~ (fsm_output[7])));
  assign mux_1185_nl = MUX_s_1_2_2((mux_1184_nl), (nor_587_nl), fsm_output[4]);
  assign nor_588_nl = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[0]) | (fsm_output[1])
      | (fsm_output[6]) | (~ (fsm_output[7])));
  assign mux_1186_nl = MUX_s_1_2_2((mux_1185_nl), (nor_588_nl), fsm_output[3]);
  assign and_658_nl = and_dcpl_624 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_447_m1c;
  assign and_659_nl = and_dcpl_626 & nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_447_m1c;
  assign or_1788_nl = (fsm_output[2]) | (fsm_output[6]) | nand_198_cse;
  assign mux_1189_nl = MUX_s_1_2_2((or_1788_nl), or_tmp_1115, fsm_output[1]);
  assign or_1786_nl = (~ (fsm_output[2])) | (~ (fsm_output[6])) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1187_nl = MUX_s_1_2_2((or_1786_nl), or_tmp_1115, fsm_output[1]);
  assign nand_177_nl = ~(IndexLoop_stage_0_2 & (~ (mux_1187_nl)));
  assign or_1784_nl = (~ (fsm_output[1])) | (fsm_output[2]) | (fsm_output[6]) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1188_nl = MUX_s_1_2_2((nand_177_nl), (or_1784_nl), IndexLoop_stage_0);
  assign mux_1190_nl = MUX_s_1_2_2((mux_1189_nl), (mux_1188_nl), fsm_output[0]);
  assign or_1783_nl = and_2642_cse | (fsm_output[6]) | nand_198_cse;
  assign mux_1191_nl = MUX_s_1_2_2((mux_1190_nl), (or_1783_nl), fsm_output[4]);
  assign or_1792_nl = (fsm_output[4]) | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1192_nl = MUX_s_1_2_2(nand_198_cse, (or_1792_nl), fsm_output[1]);
  assign nand_178_nl = ~((fsm_output[1]) & (~((~ or_tmp_940) | (fsm_output[4]) |
      (fsm_output[3]) | (fsm_output[7]))));
  assign mux_1193_nl = MUX_s_1_2_2((mux_1192_nl), (nand_178_nl), fsm_output[0]);
  assign nor_578_nl = ~((fsm_output[2]) | (mux_1193_nl));
  assign nor_580_nl = ~((fsm_output[2:0]!=3'b101) | IndexLoop_stage_0 | (~ IndexLoop_stage_0_2)
      | (fsm_output[4]) | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1194_nl = MUX_s_1_2_2((nor_578_nl), (nor_580_nl), fsm_output[6]);
  assign ReuseLoop_1_ir_ReuseLoop_1_ir_and_nl = MUX_v_11_2_2(11'b00000000000, (z_out_12[10:0]),
      and_dcpl_60);
  assign ReuseLoop_2_ir_ReuseLoop_2_ir_and_nl = MUX_v_9_2_2(9'b000000000, z_out_11,
      and_dcpl_55);
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_or_446_nl =
      and_dcpl_158 | nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_643_rgt;
  assign nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_and_845_nl
      = (~ and_dcpl_175) & and_dcpl_467;
  assign and_656_nl = and_dcpl_624 & and_dcpl_517;
  assign and_657_nl = and_dcpl_626 & and_dcpl_517;
  assign mux_949_nl = MUX_s_1_2_2(mux_tmp_774, mux_tmp_787, fsm_output[0]);
  assign mux_796_nl = MUX_s_1_2_2(mux_tmp_184, mux_tmp_530, and_2657_cse);
  assign and_627_nl = and_dcpl_624 & and_dcpl_587;
  assign and_629_nl = and_dcpl_626 & and_dcpl_587;
  assign or_1797_nl = (fsm_output[2:0]!=3'b000);
  assign mux_1197_nl = MUX_s_1_2_2(nand_tmp_65, (or_1797_nl), fsm_output[5]);
  assign or_1794_nl = (fsm_output[6]) | (fsm_output[2]) | (fsm_output[0]) | (fsm_output[1]);
  assign mux_1196_nl = MUX_s_1_2_2(nand_tmp_65, (or_1794_nl), fsm_output[5]);
  assign mux_1198_nl = MUX_s_1_2_2((mux_1197_nl), (mux_1196_nl), z_out_23_22_8[10]);
  assign and_654_nl = and_dcpl_624 & and_dcpl_579;
  assign and_655_nl = and_dcpl_626 & and_dcpl_579;
  assign mux_807_nl = MUX_s_1_2_2(mux_tmp_806, mux_tmp_742, or_1875_cse);
  assign and_630_nl = and_dcpl_624 & and_dcpl_592;
  assign and_631_nl = and_dcpl_626 & and_dcpl_592;
  assign or_1803_nl = (fsm_output[1]) | (~ (fsm_output[5])) | (fsm_output[2]);
  assign mux_1203_nl = MUX_s_1_2_2(nand_152_cse, (fsm_output[2]), fsm_output[5]);
  assign or_1802_nl = (~ (fsm_output[5])) | (fsm_output[2]);
  assign mux_1204_nl = MUX_s_1_2_2((mux_1203_nl), (or_1802_nl), IndexLoop_stage_0);
  assign mux_1205_nl = MUX_s_1_2_2((mux_1204_nl), or_tmp_1128, fsm_output[1]);
  assign mux_1206_nl = MUX_s_1_2_2((or_1803_nl), (mux_1205_nl), IndexLoop_stage_0_2);
  assign or_1801_nl = (fsm_output[1]) | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[2]);
  assign mux_1199_nl = MUX_s_1_2_2(nand_152_cse, or_1800_cse, fsm_output[5]);
  assign or_1799_nl = (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[2]);
  assign mux_1200_nl = MUX_s_1_2_2((mux_1199_nl), (or_1799_nl), IndexLoop_stage_0);
  assign mux_1201_nl = MUX_s_1_2_2((mux_1200_nl), or_tmp_1128, fsm_output[1]);
  assign mux_1202_nl = MUX_s_1_2_2((or_1801_nl), (mux_1201_nl), IndexLoop_stage_0_2);
  assign mux_1207_nl = MUX_s_1_2_2((mux_1206_nl), (mux_1202_nl), z_out_23_22_8[10]);
  assign and_652_nl = and_dcpl_624 & and_dcpl_576;
  assign and_653_nl = and_dcpl_626 & and_dcpl_576;
  assign mux_948_nl = MUX_s_1_2_2(mux_tmp_787, mux_tmp_831, fsm_output[0]);
  assign mux_821_nl = MUX_s_1_2_2(mux_tmp_806, mux_tmp_742, fsm_output[1]);
  assign mux_822_nl = MUX_s_1_2_2((mux_821_nl), mux_tmp_820, fsm_output[0]);
  assign and_632_nl = and_dcpl_624 & and_dcpl_154;
  assign and_633_nl = and_dcpl_626 & and_dcpl_154;
  assign or_1809_nl = (~ (fsm_output[5])) | (~ (fsm_output[1])) | (fsm_output[2]);
  assign mux_1211_nl = MUX_s_1_2_2((or_1809_nl), nand_tmp_66, fsm_output[0]);
  assign or_1808_nl = (~ (fsm_output[5])) | (fsm_output[6]) | (~ (fsm_output[1]))
      | (fsm_output[2]);
  assign mux_1210_nl = MUX_s_1_2_2((or_1808_nl), nand_tmp_66, fsm_output[0]);
  assign mux_1212_nl = MUX_s_1_2_2((mux_1211_nl), (mux_1210_nl), z_out_23_22_8[10]);
  assign and_650_nl = and_dcpl_624 & and_dcpl_573;
  assign and_651_nl = and_dcpl_626 & and_dcpl_573;
  assign mux_838_nl = MUX_s_1_2_2(mux_tmp_837, mux_tmp_820, fsm_output[0]);
  assign and_634_nl = and_dcpl_624 & and_dcpl_62;
  assign and_635_nl = and_dcpl_626 & and_dcpl_62;
  assign mux_1216_nl = MUX_s_1_2_2(nand_tmp_67, or_1286_cse, fsm_output[5]);
  assign mux_1215_nl = MUX_s_1_2_2(nand_tmp_67, or_tmp_1140, fsm_output[5]);
  assign mux_1217_nl = MUX_s_1_2_2((mux_1216_nl), (mux_1215_nl), z_out_23_22_8[10]);
  assign and_648_nl = and_dcpl_624 & and_dcpl_570;
  assign and_649_nl = and_dcpl_626 & and_dcpl_570;
  assign mux_947_nl = MUX_s_1_2_2(mux_tmp_831, mux_tmp_845, fsm_output[0]);
  assign and_636_nl = and_dcpl_624 & and_dcpl_157;
  assign and_637_nl = and_dcpl_626 & and_dcpl_157;
  assign mux_944_nl = MUX_s_1_2_2(mux_tmp_861, mux_tmp_837, fsm_output[0]);
  assign and_646_nl = and_dcpl_624 & and_dcpl_567;
  assign and_647_nl = and_dcpl_626 & and_dcpl_567;
  assign and_640_nl = and_dcpl_624 & and_dcpl_159;
  assign and_641_nl = and_dcpl_626 & and_dcpl_159;
  assign mux_945_nl = MUX_s_1_2_2(mux_tmp_870, mux_tmp_861, fsm_output[0]);
  assign and_644_nl = and_dcpl_624 & and_dcpl_519;
  assign and_645_nl = and_dcpl_626 & and_dcpl_519;
  assign mux_946_nl = MUX_s_1_2_2(mux_tmp_845, mux_tmp_870, fsm_output[0]);
  assign and_642_nl = and_dcpl_624 & and_dcpl_51;
  assign and_643_nl = and_dcpl_626 & and_dcpl_51;
  assign nand_183_nl = ~(IndexLoop_stage_0_2 & (~ mux_tmp_1216));
  assign or_1820_nl = (fsm_output[7]) | (fsm_output[3]) | mux_tmp_1215;
  assign mux_1221_nl = MUX_s_1_2_2(mux_tmp_1216, (or_1820_nl), and_2630_cse);
  assign mux_1222_nl = MUX_s_1_2_2((nand_183_nl), (mux_1221_nl), IndexLoop_stage_0);
  assign nor_569_nl = ~((fsm_output[6]) | (~(or_1875_cse & (fsm_output[2]))));
  assign nor_570_nl = ~((fsm_output[6]) | and_2642_cse);
  assign mux_1218_nl = MUX_s_1_2_2((nor_569_nl), (nor_570_nl), fsm_output[3]);
  assign nand_182_nl = ~((fsm_output[7]) & (mux_1218_nl));
  assign mux_1223_nl = MUX_s_1_2_2((mux_1222_nl), (nand_182_nl), fsm_output[4]);
  assign nor_571_nl = ~((~ (fsm_output[1])) | (fsm_output[6]) | (fsm_output[7]) |
      or_1876_cse);
  assign nor_572_nl = ~((fsm_output[7]) | or_1876_cse);
  assign mux_1225_nl = MUX_s_1_2_2(and_2631_cse, (nor_572_nl), fsm_output[6]);
  assign or_1825_nl = IndexLoop_stage_0 | (~ IndexLoop_stage_0_2) | (fsm_output[4]);
  assign mux_1224_nl = MUX_s_1_2_2(or_1876_cse, (or_1825_nl), and_2630_cse);
  assign nor_573_nl = ~((fsm_output[7:6]!=2'b10) | (mux_1224_nl));
  assign mux_1226_nl = MUX_s_1_2_2((mux_1225_nl), (nor_573_nl), fsm_output[1]);
  assign mux_1227_nl = MUX_s_1_2_2((nor_571_nl), (mux_1226_nl), fsm_output[2]);
  assign and_2625_nl = (fsm_output[4]) & (fsm_output[7]) & (fsm_output[3]);
  assign nor_558_nl = ~((fsm_output[4]) | (fsm_output[7]) | (~(or_tmp_940 & (fsm_output[0])
      & (fsm_output[2]) & (~ (fsm_output[3])))));
  assign mux_1234_nl = MUX_s_1_2_2((and_2625_nl), (nor_558_nl), fsm_output[6]);
  assign or_1837_nl = ((~((~(nand_191_cse & IndexLoop_stage_0)) & IndexLoop_stage_0_2))
      & (fsm_output[0])) | (fsm_output[3:2]!=2'b00);
  assign nand_192_nl = ~(IndexLoop_stage_0_2 & (fsm_output[0]) & (fsm_output[2])
      & (~ (fsm_output[3])));
  assign or_1834_nl = (MultLoop_2_1_acc_3_tmp[1]) | (~ (fsm_output[0])) | (~ (fsm_output[2]))
      | (fsm_output[3]);
  assign or_1833_nl = nor_560_cse | (~ (fsm_output[0])) | (~ (fsm_output[2])) | (fsm_output[3]);
  assign mux_1230_nl = MUX_s_1_2_2((or_1834_nl), (or_1833_nl), MultLoop_2_1_acc_3_tmp[2]);
  assign mux_1231_nl = MUX_s_1_2_2((nand_192_nl), (mux_1230_nl), IndexLoop_stage_0);
  assign mux_1232_nl = MUX_s_1_2_2((or_1837_nl), (mux_1231_nl), fsm_output[7]);
  assign mux_1228_nl = MUX_s_1_2_2((fsm_output[3]), (~ (fsm_output[3])), fsm_output[2]);
  assign mux_1229_nl = MUX_s_1_2_2(or_647_cse_1, (mux_1228_nl), fsm_output[0]);
  assign nand_185_nl = ~((fsm_output[7]) & (mux_1229_nl));
  assign mux_1233_nl = MUX_s_1_2_2((mux_1232_nl), (nand_185_nl), fsm_output[4]);
  assign nor_559_nl = ~((fsm_output[6]) | (mux_1233_nl));
  assign mux_1235_nl = MUX_s_1_2_2((mux_1234_nl), (nor_559_nl), fsm_output[1]);
  assign nor_561_nl = ~((fsm_output[2]) | (fsm_output[4]));
  assign and_2628_nl = (fsm_output[2]) & (fsm_output[4]);
  assign mux_1239_nl = MUX_s_1_2_2((nor_561_nl), (and_2628_nl), fsm_output[7]);
  assign nor_562_nl = ~((nand_191_cse & IndexLoop_stage_0) | (~ IndexLoop_stage_0_2)
      | (fsm_output[2]) | (fsm_output[4]));
  assign nor_563_nl = ~((~ IndexLoop_stage_0_2) | (~ (fsm_output[2])) | (fsm_output[4]));
  assign nor_564_nl = ~((MultLoop_2_1_acc_3_tmp[1]) | (~ (fsm_output[2])) | (fsm_output[4]));
  assign nor_565_nl = ~(nor_560_cse | (~ (fsm_output[2])) | (fsm_output[4]));
  assign mux_1236_nl = MUX_s_1_2_2((nor_564_nl), (nor_565_nl), MultLoop_2_1_acc_3_tmp[2]);
  assign mux_1237_nl = MUX_s_1_2_2((nor_563_nl), (mux_1236_nl), IndexLoop_stage_0);
  assign mux_1238_nl = MUX_s_1_2_2((nor_562_nl), (mux_1237_nl), fsm_output[7]);
  assign mux_1240_nl = MUX_s_1_2_2((mux_1239_nl), (mux_1238_nl), fsm_output[0]);
  assign and_2627_nl = (fsm_output[1]) & (mux_1240_nl);
  assign nor_567_nl = ~((fsm_output[1]) | (~ (fsm_output[0])) | (fsm_output[7]) |
      (~ or_tmp_940) | (~ (fsm_output[2])) | (fsm_output[4]));
  assign mux_1241_nl = MUX_s_1_2_2((and_2627_nl), (nor_567_nl), fsm_output[6]);
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_194_nl
      = (and_dcpl_424 & and_dcpl_261 & and_dcpl_65) | ((~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_126_tmp)
      & and_dcpl_60);
  assign MultLoop_and_215_nl = (~ or_dcpl_588) & and_554_m1c & and_dcpl_65;
  assign MultLoop_and_216_nl = or_dcpl_588 & and_554_m1c & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_and_136_nl
      = (~ or_dcpl_490) & and_dcpl_158;
  assign and_555_nl = and_dcpl_326 & and_dcpl_261 & and_dcpl_65;
  assign nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_195_nl
      = ((~ or_dcpl_590) & and_556_m1c & and_dcpl_65) | ((~ nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_or_127_tmp)
      & and_dcpl_60);
  assign MultLoop_and_212_nl = or_dcpl_590 & and_556_m1c & and_dcpl_65;
  assign and_557_nl = and_dcpl_64 & and_dcpl_159;
  assign and_560_nl = ((and_817_cse & (fsm_output[0])) ^ (fsm_output[3])) & and_dcpl_100;
  assign and_562_nl = and_dcpl_54 & and_dcpl_57;
  assign or_1358_nl = (or_1405_cse & (fsm_output[6])) | (fsm_output[7]);
  assign mux_916_nl = MUX_s_1_2_2(mux_tmp_914, (or_1358_nl), fsm_output[2]);
  assign mux_917_nl = MUX_s_1_2_2((mux_916_nl), mux_tmp_915, fsm_output[1]);
  assign mux_919_nl = MUX_s_1_2_2(mux_tmp_918, (mux_917_nl), fsm_output[0]);
  assign and_564_nl = and_dcpl_54 & and_dcpl_157;
  assign mux_920_nl = MUX_s_1_2_2(mux_661_cse, or_tmp_91, or_1405_cse);
  assign mux_921_nl = MUX_s_1_2_2(mux_tmp_914, (mux_920_nl), fsm_output[2]);
  assign mux_922_nl = MUX_s_1_2_2((mux_921_nl), mux_tmp_915, fsm_output[1]);
  assign mux_923_nl = MUX_s_1_2_2(mux_tmp_918, (mux_922_nl), fsm_output[0]);
  assign and_571_nl = and_dcpl_59 & and_dcpl_567;
  assign and_574_nl = and_dcpl_59 & and_dcpl_570;
  assign mux_929_nl = MUX_s_1_2_2(mux_tmp_928, mux_tmp_926, fsm_output[0]);
  assign and_577_nl = and_dcpl_59 & and_dcpl_573;
  assign and_580_nl = and_dcpl_59 & and_dcpl_576;
  assign mux_931_nl = MUX_s_1_2_2(mux_tmp_930, mux_tmp_928, fsm_output[0]);
  assign and_583_nl = and_dcpl_59 & and_dcpl_579;
  assign and_585_nl = and_dcpl_59 & and_dcpl_517;
  assign mux_932_nl = MUX_s_1_2_2(mux_tmp_500, mux_tmp_930, fsm_output[0]);
  assign and_610_nl = and_dcpl_590 & and_dcpl_519;
  assign mux_938_nl = MUX_s_1_2_2(mux_tmp_707, mux_tmp_670, fsm_output[0]);
  assign and_624_nl = and_dcpl_590 & and_dcpl_584;
  assign mux_800_nl = MUX_s_1_2_2(mux_tmp_184, mux_tmp_530, and_817_cse);
  assign or_1868_nl = (fsm_output[4:3]!=2'b10);
  assign or_1867_nl = (fsm_output[4:3]!=2'b01);
  assign mux_1247_nl = MUX_s_1_2_2((or_1868_nl), (or_1867_nl), fsm_output[2]);
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_nor_nl
      = ~((z_out_10!=71'b00000000000000000000000000000000000000000000000000000000000000000000000));
  assign ReuseLoop_1_ReuseLoop_1_mux_1_nl = MUX_v_6_2_2(InitAccumLoop_1_iacc_6_0_sva_5_0,
      ({5'b00000 , (~ (IndexLoop_if_acc_3_psp_1_sva_1[5]))}), and_dcpl_737);
  assign ReuseLoop_1_or_3_nl = (~(and_dcpl_730 | and_dcpl_741)) | and_dcpl_737;
  assign ReuseLoop_1_or_4_nl = (IndexLoop_if_acc_3_psp_1_sva_1[6]) | and_dcpl_730
      | and_dcpl_741;
  assign nl_acc_nl = conv_u2u_7_8({(ReuseLoop_1_ReuseLoop_1_mux_1_nl) , (ReuseLoop_1_or_3_nl)})
      + conv_u2u_2_8({(ReuseLoop_1_or_4_nl) , 1'b1});
  assign acc_nl = nl_acc_nl[7:0];
  assign z_out = readslicef_8_7_1((acc_nl));
  assign and_2668_nl = (fsm_output[7:6]==2'b10) & (~((fsm_output[4]) ^ (fsm_output[3])))
      & (~ (fsm_output[5])) & (fsm_output[2]) & (fsm_output[1]) & (~ (fsm_output[0]));
  assign ReuseLoop_2_mux_1_nl = MUX_v_3_2_2((z_out_11[8:6]), (z_out_4[3:1]), and_2668_nl);
  assign nl_ReuseLoop_2_acc_nl = conv_u2u_3_4(ReuseLoop_2_mux_1_nl) + 4'b1011;
  assign ReuseLoop_2_acc_nl = nl_ReuseLoop_2_acc_nl[3:0];
  assign z_out_1_3 = readslicef_4_1_3((ReuseLoop_2_acc_nl));
  assign ac_math_ac_reciprocal_pwl_AC_TRN_71_51_false_AC_TRN_AC_WRAP_91_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_71_51_false_AC_TRN_AC_WRAP_91_21_false_AC_TRN_AC_WRAP_output_pwl_or_1_nl
      = (~(and_dcpl_764 | and_dcpl_768)) | and_dcpl_760;
  assign ac_math_ac_reciprocal_pwl_AC_TRN_71_51_false_AC_TRN_AC_WRAP_91_21_false_AC_TRN_AC_WRAP_output_pwl_mux1h_2_nl
      = MUX1HOT_v_10_3_2(ROM_1i3_1o10_bb905e8578f158e8f5b59add1dc96bdb2f_1, reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd_2,
      10'b0000000101, {and_dcpl_760 , and_dcpl_764 , and_dcpl_768});
  assign ac_math_ac_reciprocal_pwl_AC_TRN_71_51_false_AC_TRN_AC_WRAP_91_21_false_AC_TRN_AC_WRAP_output_pwl_mux1h_3_nl
      = MUX1HOT_v_9_3_2((z_out_17[18:10]), 9'b000000001, ({6'b000000 , (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2[8:6])}),
      {and_dcpl_760 , and_dcpl_764 , and_dcpl_768});
  assign nl_z_out_2 = ({(ac_math_ac_reciprocal_pwl_AC_TRN_71_51_false_AC_TRN_AC_WRAP_91_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_71_51_false_AC_TRN_AC_WRAP_91_21_false_AC_TRN_AC_WRAP_output_pwl_or_1_nl)
      , (ac_math_ac_reciprocal_pwl_AC_TRN_71_51_false_AC_TRN_AC_WRAP_91_21_false_AC_TRN_AC_WRAP_output_pwl_mux1h_2_nl)})
      + conv_s2u_9_11(ac_math_ac_reciprocal_pwl_AC_TRN_71_51_false_AC_TRN_AC_WRAP_91_21_false_AC_TRN_AC_WRAP_output_pwl_mux1h_3_nl);
  assign z_out_2 = nl_z_out_2[10:0];
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_qif_mux_2_nl = MUX_v_6_2_2(({1'b1
      , (~ (libraries_leading_sign_71_0_e5d4bd9dc928fda5adf5bf26ec9a2550b9a2_1[6:2]))}),
      (IndexLoop_if_acc_4_psp_sva_1[5:0]), and_dcpl_779);
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_qif_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_qif_and_1_nl
      = (IndexLoop_if_acc_4_psp_sva_1[6]) & and_dcpl_779;
  assign ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_qif_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_qif_or_1_nl
      = (IndexLoop_if_acc_4_psp_sva_1[6]) | (~ and_dcpl_779);
  assign nl_z_out_3 = (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_qif_mux_2_nl)
      + conv_s2u_5_6({(ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_qif_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_qif_and_1_nl)
      , (~ and_dcpl_779) , (~ and_dcpl_779) , 1'b0 , (ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_qif_ac_math_ac_normalize_71_51_false_AC_TRN_AC_WRAP_expret_qif_or_1_nl)});
  assign z_out_3 = nl_z_out_3[5:0];
  assign nl_z_out_4 = InitAccumLoop_2_iacc_3_0_sva + 4'b0001;
  assign z_out_4 = nl_z_out_4[3:0];
  assign SUM_EXP_LOOP_SUM_EXP_LOOP_and_5_nl = (SUM_EXP_LOOP_acc_itm_69_68[1]) & SUM_EXP_LOOP_nor_itm;
  assign SUM_EXP_LOOP_mux_3_nl = MUX_s_1_2_2((z_out_24[68]), (SUM_EXP_LOOP_acc_itm_69_68[0]),
      and_dcpl_967);
  assign SUM_EXP_LOOP_SUM_EXP_LOOP_and_6_nl = (SUM_EXP_LOOP_mux_3_nl) & (~ and_dcpl_964);
  assign SUM_EXP_LOOP_or_1_nl = and_dcpl_964 | and_dcpl_967;
  assign SUM_EXP_LOOP_SUM_EXP_LOOP_mux_2_nl = MUX_v_68_2_2((z_out_24[67:0]), SUM_EXP_LOOP_acc_itm_67_0,
      SUM_EXP_LOOP_or_1_nl);
  assign SUM_EXP_LOOP_SUM_EXP_LOOP_and_7_nl = (SUM_EXP_LOOP_acc_11_itm[68]) & SUM_EXP_LOOP_nor_itm;
  assign SUM_EXP_LOOP_mux1h_5_nl = MUX1HOT_v_68_3_2(SUM_EXP_LOOP_acc_9_itm, (z_out_24[67:0]),
      (SUM_EXP_LOOP_acc_11_itm[67:0]), {and_1134_cse , and_dcpl_964 , and_dcpl_967});
  assign nl_z_out_10 = conv_u2u_70_71({(SUM_EXP_LOOP_SUM_EXP_LOOP_and_5_nl) , (SUM_EXP_LOOP_SUM_EXP_LOOP_and_6_nl)
      , (SUM_EXP_LOOP_SUM_EXP_LOOP_mux_2_nl)}) + conv_u2u_69_71({(SUM_EXP_LOOP_SUM_EXP_LOOP_and_7_nl)
      , (SUM_EXP_LOOP_mux1h_5_nl)});
  assign z_out_10 = nl_z_out_10[70:0];
  assign ReuseLoop_if_mux_2_nl = MUX_v_9_2_2(({2'b00 , (z_out_2[10:4])}), (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2[8:0]),
      and_dcpl_979);
  assign nl_z_out_11 = (ReuseLoop_if_mux_2_nl) + conv_s2u_7_9({(~ and_dcpl_979) ,
      2'b00 , (signext_3_1(~ and_dcpl_979)) , 1'b1});
  assign z_out_11 = nl_z_out_11[8:0];
  assign ReuseLoop_mux1h_5_nl = MUX1HOT_s_1_10_2((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg[2]),
      (reg_MultLoop_1_mux_64_itm_1_reg[5]), (reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_reg[5]),
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_1_ftd,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_1_ftd,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_1_ftd,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd,
      (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2[17]),
      {and_1173_cse , and_1175_cse , and_1178_cse , and_1180_cse , and_1183_cse ,
      and_1185_cse , and_1187_cse , and_1189_cse , and_1193_cse , and_1195_cse});
  assign ReuseLoop_and_4_nl = (ReuseLoop_mux1h_5_nl) & ReuseLoop_nor_itm;
  assign ReuseLoop_mux1h_6_nl = MUX1HOT_v_15_10_2(nnet_softmax_layer6_t_result_t_softmax_config7_for_1_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_psp_sva_1,
      ({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_2_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_4_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2}),
      ({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_1_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_2_reg}),
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_14_0,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_14_0,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_14_0,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_14_0,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_14_0,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_14_0,
      ({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_2_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg}),
      {and_1173_cse , and_1175_cse , and_1178_cse , and_1180_cse , and_1183_cse ,
      and_1185_cse , and_1187_cse , and_1189_cse , and_1193_cse , and_1195_cse});
  assign ReuseLoop_and_5_nl = MUX_v_15_2_2(15'b000000000000000, (ReuseLoop_mux1h_6_nl),
      ReuseLoop_nor_itm);
  assign ReuseLoop_mux_1_nl = MUX_v_8_2_2((signext_8_4({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_2_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_4_reg})),
      (z_out_13[21:14]), ReuseLoop_or_itm);
  assign not_3912_nl = ~ and_dcpl_992;
  assign ReuseLoop_ReuseLoop_and_2_nl = MUX_v_8_2_2(8'b00000000, (ReuseLoop_mux_1_nl),
      (not_3912_nl));
  assign ReuseLoop_ReuseLoop_mux_1_nl = MUX_v_11_2_2(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2,
      (z_out_13[13:3]), ReuseLoop_or_itm);
  assign nl_z_out_12 = ({(ReuseLoop_and_4_nl) , (ReuseLoop_and_5_nl) , ReuseLoop_and_2_cse
      , ReuseLoop_and_2_cse , 2'b01}) + conv_s2u_19_20({(ReuseLoop_ReuseLoop_and_2_nl)
      , (ReuseLoop_ReuseLoop_mux_1_nl)});
  assign z_out_12 = nl_z_out_12[19:0];
  assign IndexLoop_if_mux1h_5_nl = MUX1HOT_s_1_11_2((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_2_reg[2]),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg[2])),
      (~ (reg_MultLoop_1_mux_64_itm_1_reg[5])), (~ (reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_reg[5])),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd),
      (~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2[17])),
      {and_1161_cse , and_1173_cse , and_1175_cse , and_1178_cse , and_1180_cse ,
      and_1183_cse , and_1185_cse , and_1187_cse , and_1189_cse , and_1193_cse ,
      and_1195_cse});
  assign IndexLoop_if_mux1h_6_nl = MUX1HOT_v_15_11_2((signext_15_10({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_2_reg
      , (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg[11:5])})),
      (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_1_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_psp_sva_1),
      ({(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_2_reg)
      , (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_4_reg)
      , (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2)}),
      ({(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_1_reg)
      , (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_2_reg)}),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_14_0),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_14_0),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_14_0),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_14_0),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_14_0),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_14_0),
      ({(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_2_reg)
      , (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg)}),
      {and_1161_cse , and_1173_cse , and_1175_cse , and_1178_cse , and_1180_cse ,
      and_1183_cse , and_1185_cse , and_1187_cse , and_1189_cse , and_1193_cse ,
      and_1195_cse});
  assign IndexLoop_if_mux1h_7_nl = MUX1HOT_s_1_11_2((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg[4]),
      (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_1_sva_1), (~
      MultLoop_2_and_5_itm_1), (~ MultLoop_2_and_6_itm_1), (~ MultLoop_2_and_7_itm_1),
      (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_5_sva), (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_6_sva),
      (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_7_sva), (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_8_sva),
      (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_9_sva), (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_sva),
      {and_1161_cse , and_1173_cse , and_1175_cse , and_1178_cse , and_1180_cse ,
      and_1183_cse , and_1185_cse , and_1187_cse , and_1189_cse , and_1193_cse ,
      and_1195_cse});
  assign IndexLoop_if_mux1h_8_nl = MUX1HOT_s_1_11_2((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg[3]),
      (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_1_sva_1), (~
      MultLoop_2_and_5_itm_1), (~ MultLoop_2_and_6_itm_1), (~ MultLoop_2_and_7_itm_1),
      (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_5_sva), (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_6_sva),
      (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_7_sva), (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_8_sva),
      (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_9_sva), (~ nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_sva),
      {and_1161_cse , and_1173_cse , and_1175_cse , and_1178_cse , and_1180_cse ,
      and_1183_cse , and_1185_cse , and_1187_cse , and_1189_cse , and_1193_cse ,
      and_1195_cse});
  assign IndexLoop_if_IndexLoop_if_and_2_nl = (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg[2])
      & IndexLoop_if_nor_itm;
  assign IndexLoop_if_IndexLoop_if_and_3_nl = (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg[1])
      & IndexLoop_if_nor_itm;
  assign IndexLoop_if_IndexLoop_if_or_1_nl = (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg[0])
      | and_1173_cse | and_1175_cse | and_1178_cse | and_1180_cse | and_1183_cse
      | and_1185_cse | and_1187_cse | and_1189_cse | and_1193_cse | and_1195_cse;
  assign ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_17_nl
      = MUX1HOT_s_1_10_2((~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg[2])),
      (~ (reg_MultLoop_1_mux_64_itm_1_reg[5])), (~ (reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_reg[5])),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd),
      (~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2[17])),
      {and_1270_cse , and_1273_cse , and_1276_cse , and_1279_cse , and_1282_cse ,
      and_1284_cse , and_1286_cse , and_1288_cse , and_1193_cse , and_1195_cse});
  assign ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_18_nl
      = MUX1HOT_v_15_10_2((~ nnet_softmax_layer6_t_result_t_softmax_config7_for_1_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_psp_sva_1),
      ({(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_2_reg)
      , (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_4_reg)
      , (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2)}),
      ({(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_1_reg)
      , (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_2_reg)}),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_14_0),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_14_0),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_14_0),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_14_0),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_14_0),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_14_0),
      ({(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_2_reg)
      , (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg)}),
      {and_1270_cse , and_1273_cse , and_1276_cse , and_1279_cse , and_1282_cse ,
      and_1284_cse , and_1286_cse , and_1288_cse , and_1193_cse , and_1195_cse});
  assign nl_ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_80_nl
      = ({(ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_17_nl)
      , (ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_18_nl)
      , ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_7_cse
      , ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_7_cse})
      + conv_s2u_15_18(z_out_23_22_8);
  assign ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_80_nl
      = nl_ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_80_nl[17:0];
  assign IndexLoop_if_IndexLoop_if_mux_1_nl = MUX_v_18_2_2(18'b000000000000000001,
      (ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_80_nl),
      ReuseLoop_or_itm);
  assign nl_z_out_13 = conv_s2u_21_22({(IndexLoop_if_mux1h_5_nl) , (IndexLoop_if_mux1h_6_nl)
      , (IndexLoop_if_mux1h_7_nl) , (IndexLoop_if_mux1h_8_nl) , (IndexLoop_if_IndexLoop_if_and_2_nl)
      , (IndexLoop_if_IndexLoop_if_and_3_nl) , (IndexLoop_if_IndexLoop_if_or_1_nl)})
      + conv_s2u_18_22(IndexLoop_if_IndexLoop_if_mux_1_nl);
  assign z_out_13 = nl_z_out_13[21:0];
  assign ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_19_cse
      = MUX1HOT_v_15_10_2(nnet_softmax_layer6_t_result_t_softmax_config7_for_1_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_psp_sva_1,
      ({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_2_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_4_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2}),
      ({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_1_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_2_reg}),
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_14_0,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_14_0,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_14_0,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_14_0,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_14_0,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_14_0,
      ({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_2_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg}),
      {and_1270_cse , and_1273_cse , and_1276_cse , and_1279_cse , and_1282_cse ,
      and_1284_cse , and_1286_cse , and_1288_cse , and_1193_cse , and_1195_cse});
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_mux_2_nl = MUX_v_18_2_2(MultLoop_1_slc_input1_18_17_0_cse_sva_1,
      ({10'b1111111111 , ROM_1i3_1o8_bdb5a3eca137308489a677a1241b230a2e_1}), and_dcpl_1163);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_mux_3_nl = MUX_v_18_2_2((w2_rsci_qa_d_mxwt[17:0]),
      ({8'b00000000 , (operator_71_0_false_AC_TRN_AC_WRAP_lshift_itm[66:57])}), and_dcpl_1163);
  assign nl_z_out_17 = $signed((nnet_product_input_t_config2_weight_t_config2_accum_t_mux_2_nl))
      * $signed((nnet_product_input_t_config2_weight_t_config2_accum_t_mux_3_nl));
  assign z_out_17 = nl_z_out_17[27:0];
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_1_or_2_nl = and_dcpl_1170
      | and_dcpl_1175;
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_1_mux1h_3_nl = MUX1HOT_v_67_11_2(({50'b00000000000000000000000000000000000000000000000000
      , (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_1_ftd[1:0])
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_2_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg}),
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_10_18_6_true_AC_TRN_AC_SAT_18_2_AC_TRN_AC_SAT_exp_arr_0_sva,
      CALC_EXP_LOOP_2_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva, CALC_EXP_LOOP_3_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva,
      CALC_EXP_LOOP_4_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva, CALC_EXP_LOOP_5_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva,
      CALC_EXP_LOOP_6_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva, CALC_EXP_LOOP_7_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva,
      CALC_EXP_LOOP_8_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva, CALC_EXP_LOOP_9_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva,
      CALC_EXP_LOOP_10_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva, {(nnet_product_input_t_config2_weight_t_config2_accum_t_1_or_2_nl)
      , and_dcpl_1180 , and_dcpl_1181 , and_dcpl_1184 , and_dcpl_1185 , and_dcpl_1188
      , and_dcpl_1190 , and_dcpl_1192 , and_dcpl_1194 , and_dcpl_1197 , and_dcpl_1199});
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_1_mux_3_nl = MUX_s_1_2_2((w4_rsci_qa_d_mxwt[35]),
      (w6_rsci_qa_d_mxwt[35]), and_dcpl_1175);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_1_nnet_product_input_t_config2_weight_t_config2_accum_t_1_and_1_nl
      = (nnet_product_input_t_config2_weight_t_config2_accum_t_1_mux_3_nl) & (~(and_dcpl_1180
      | and_dcpl_1181 | and_dcpl_1184 | and_dcpl_1185 | and_dcpl_1188 | and_dcpl_1190
      | and_dcpl_1192 | and_dcpl_1194 | and_dcpl_1197 | and_dcpl_1199));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_1_mux1h_4_nl = MUX1HOT_v_74_3_2((signext_74_1(w4_rsci_qa_d_mxwt[35])),
      (signext_74_1(w6_rsci_qa_d_mxwt[35])), (ac_math_ac_reciprocal_pwl_AC_TRN_71_51_false_AC_TRN_AC_WRAP_91_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1_dfm[90:17]),
      {and_dcpl_1170 , and_dcpl_1175 , nnet_product_input_t_config2_weight_t_config2_accum_t_1_or_1_ssc});
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_1_mux1h_5_nl = MUX1HOT_v_17_3_2((w4_rsci_qa_d_mxwt[34:18]),
      (w6_rsci_qa_d_mxwt[34:18]), (ac_math_ac_reciprocal_pwl_AC_TRN_71_51_false_AC_TRN_AC_WRAP_91_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1_dfm[16:0]),
      {and_dcpl_1170 , and_dcpl_1175 , nnet_product_input_t_config2_weight_t_config2_accum_t_1_or_1_ssc});
  assign nl_mul_1_nl = $signed(conv_u2s_67_68(nnet_product_input_t_config2_weight_t_config2_accum_t_1_mux1h_3_nl))
      * $signed(({(nnet_product_input_t_config2_weight_t_config2_accum_t_1_nnet_product_input_t_config2_weight_t_config2_accum_t_1_and_1_nl)
      , (nnet_product_input_t_config2_weight_t_config2_accum_t_1_mux1h_4_nl) , (nnet_product_input_t_config2_weight_t_config2_accum_t_1_mux1h_5_nl)}));
  assign mul_1_nl = nl_mul_1_nl[157:0];
  assign z_out_18_157_10 = readslicef_158_148_10((mul_1_nl));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_1_mux_4_nl = MUX_v_18_2_2((w4_rsci_qa_d_mxwt[17:0]),
      (w6_rsci_qa_d_mxwt[17:0]), and_dcpl_979);
  assign nl_mul_2_nl = $signed(conv_u2s_17_18({(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_1_ftd[1:0])
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_2_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg}))
      * $signed((nnet_product_input_t_config2_weight_t_config2_accum_t_1_mux_4_nl));
  assign mul_2_nl = nl_mul_2_nl[27:0];
  assign z_out_19_27_10 = readslicef_28_18_10((mul_2_nl));
  assign and_2670_cse = nor_944_cse & nor_943_cse & nor_942_cse & and_810_cse_1;
  assign MultLoop_mux_327_nl = MUX_v_18_2_2(z_out_21, ({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_1_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_2_reg}),
      or_dcpl_490);
  assign MultLoop_mux_328_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_1_1_sva_1,
      or_dcpl_372);
  assign MultLoop_mux_329_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_sva_1,
      or_dcpl_382);
  assign MultLoop_mux_330_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_sva_1,
      or_dcpl_384);
  assign MultLoop_mux_331_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_sva_1,
      or_dcpl_388);
  assign MultLoop_mux_332_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_sva_1,
      or_dcpl_390);
  assign MultLoop_mux_333_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_6_1_sva_1,
      or_dcpl_394);
  assign MultLoop_mux_334_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_sva_1,
      or_dcpl_396);
  assign MultLoop_mux_335_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_8_1_sva_1,
      or_dcpl_400);
  assign MultLoop_mux_336_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_9_1_sva_1,
      or_dcpl_404);
  assign MultLoop_mux_337_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_10_1_sva_1,
      or_dcpl_406);
  assign MultLoop_mux_338_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_sva_1,
      or_dcpl_408);
  assign MultLoop_mux_339_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_sva_1,
      or_dcpl_410);
  assign MultLoop_mux_340_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_sva_1,
      or_dcpl_412);
  assign MultLoop_mux_341_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_sva_1,
      or_dcpl_414);
  assign MultLoop_mux_342_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_sva_1,
      or_dcpl_416);
  assign MultLoop_mux_343_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_sva_1,
      or_dcpl_418);
  assign MultLoop_mux_344_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_1,
      or_dcpl_420);
  assign MultLoop_mux_345_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_sva_1,
      or_dcpl_422);
  assign MultLoop_mux_346_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_sva_1,
      or_dcpl_424);
  assign MultLoop_mux_347_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_sva_1,
      or_dcpl_426);
  assign MultLoop_mux_348_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_sva_1,
      or_dcpl_428);
  assign MultLoop_mux_349_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_sva_1,
      or_dcpl_430);
  assign MultLoop_mux_350_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_sva_1,
      or_dcpl_432);
  assign MultLoop_mux_351_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_sva_1,
      or_dcpl_434);
  assign MultLoop_mux_352_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_sva_1,
      or_dcpl_436);
  assign MultLoop_mux_353_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_sva_1,
      or_dcpl_438);
  assign MultLoop_mux_354_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_sva_1,
      or_dcpl_440);
  assign MultLoop_mux_355_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_sva_1,
      or_dcpl_442);
  assign MultLoop_mux_356_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_sva_1,
      or_dcpl_444);
  assign MultLoop_mux_357_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_sva_1,
      or_dcpl_446);
  assign MultLoop_mux_358_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_sva_1,
      or_dcpl_448);
  assign MultLoop_mux_359_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_sva_1,
      or_dcpl_447);
  assign MultLoop_mux_360_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_sva_1,
      or_dcpl_445);
  assign MultLoop_mux_361_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_sva_1,
      or_dcpl_443);
  assign MultLoop_mux_362_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_sva_1,
      or_dcpl_441);
  assign MultLoop_mux_363_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_sva_1,
      or_dcpl_439);
  assign MultLoop_mux_364_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_sva_1,
      or_dcpl_437);
  assign MultLoop_mux_365_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_sva_1,
      or_dcpl_435);
  assign MultLoop_mux_366_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_sva_1,
      or_dcpl_433);
  assign MultLoop_mux_367_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_sva_1,
      or_dcpl_431);
  assign MultLoop_mux_368_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_sva_1,
      or_dcpl_429);
  assign MultLoop_mux_369_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_sva_1,
      or_dcpl_427);
  assign MultLoop_mux_370_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_sva_1,
      or_dcpl_425);
  assign MultLoop_mux_371_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_sva_1,
      or_dcpl_423);
  assign MultLoop_mux_372_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_sva_1,
      or_dcpl_421);
  assign MultLoop_mux_373_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_sva_1,
      or_dcpl_419);
  assign MultLoop_mux_374_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_sva_1,
      or_dcpl_417);
  assign MultLoop_mux_375_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_sva_1,
      or_dcpl_415);
  assign MultLoop_mux_376_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_sva_1,
      or_dcpl_413);
  assign MultLoop_mux_377_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_sva_1,
      or_dcpl_411);
  assign MultLoop_mux_378_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_sva_1,
      or_dcpl_409);
  assign MultLoop_mux_379_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_sva_1,
      or_dcpl_407);
  assign MultLoop_mux_380_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_sva_1,
      or_dcpl_405);
  assign MultLoop_mux_381_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_sva_1,
      or_dcpl_402);
  assign MultLoop_mux_382_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_sva_1,
      or_dcpl_398);
  assign MultLoop_mux_383_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_sva_1,
      or_dcpl_395);
  assign MultLoop_mux_384_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_sva_1,
      or_dcpl_392);
  assign MultLoop_mux_385_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_58_1_sva_1,
      or_dcpl_389);
  assign MultLoop_mux_386_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_59_1_sva_1,
      or_dcpl_386);
  assign MultLoop_mux_387_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_60_1_sva_1,
      or_dcpl_383);
  assign MultLoop_mux_388_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_61_1_sva_1,
      or_dcpl_377);
  assign MultLoop_mux_389_nl = MUX_v_18_2_2(z_out_21, nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_sva_1,
      or_dcpl_366);
  assign MultLoop_mux_390_nl = MUX_v_18_2_2(z_out_21, ({reg_MultLoop_1_mux_64_itm_1_reg
      , reg_MultLoop_1_mux_64_itm_1_1_reg}), or_dcpl_560);
  assign MultLoop_mux_326_nl = MUX_v_18_64_2((MultLoop_mux_327_nl), (MultLoop_mux_328_nl),
      (MultLoop_mux_329_nl), (MultLoop_mux_330_nl), (MultLoop_mux_331_nl), (MultLoop_mux_332_nl),
      (MultLoop_mux_333_nl), (MultLoop_mux_334_nl), (MultLoop_mux_335_nl), (MultLoop_mux_336_nl),
      (MultLoop_mux_337_nl), (MultLoop_mux_338_nl), (MultLoop_mux_339_nl), (MultLoop_mux_340_nl),
      (MultLoop_mux_341_nl), (MultLoop_mux_342_nl), (MultLoop_mux_343_nl), (MultLoop_mux_344_nl),
      (MultLoop_mux_345_nl), (MultLoop_mux_346_nl), (MultLoop_mux_347_nl), (MultLoop_mux_348_nl),
      (MultLoop_mux_349_nl), (MultLoop_mux_350_nl), (MultLoop_mux_351_nl), (MultLoop_mux_352_nl),
      (MultLoop_mux_353_nl), (MultLoop_mux_354_nl), (MultLoop_mux_355_nl), (MultLoop_mux_356_nl),
      (MultLoop_mux_357_nl), (MultLoop_mux_358_nl), (MultLoop_mux_359_nl), (MultLoop_mux_360_nl),
      (MultLoop_mux_361_nl), (MultLoop_mux_362_nl), (MultLoop_mux_363_nl), (MultLoop_mux_364_nl),
      (MultLoop_mux_365_nl), (MultLoop_mux_366_nl), (MultLoop_mux_367_nl), (MultLoop_mux_368_nl),
      (MultLoop_mux_369_nl), (MultLoop_mux_370_nl), (MultLoop_mux_371_nl), (MultLoop_mux_372_nl),
      (MultLoop_mux_373_nl), (MultLoop_mux_374_nl), (MultLoop_mux_375_nl), (MultLoop_mux_376_nl),
      (MultLoop_mux_377_nl), (MultLoop_mux_378_nl), (MultLoop_mux_379_nl), (MultLoop_mux_380_nl),
      (MultLoop_mux_381_nl), (MultLoop_mux_382_nl), (MultLoop_mux_383_nl), (MultLoop_mux_384_nl),
      (MultLoop_mux_385_nl), (MultLoop_mux_386_nl), (MultLoop_mux_387_nl), (MultLoop_mux_388_nl),
      (MultLoop_mux_389_nl), (MultLoop_mux_390_nl), {(~ (InitAccumLoop_1_iacc_6_0_sva_5_0[5]))
      , (InitAccumLoop_1_iacc_6_0_sva_5_0[4:0])});
  assign MultLoop_or_9_nl = and_dcpl_1224 | and_dcpl_1228;
  assign MultLoop_mux_325_nl = MUX_v_18_2_2((MultLoop_mux_326_nl), ({reg_MultLoop_1_mux_64_itm_1_reg
      , reg_MultLoop_1_mux_64_itm_1_1_reg}), MultLoop_or_9_nl);
  assign nl_MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_1_nl
      = $signed(MultLoop_1_slc_input1_18_17_0_cse_sva_1) * $signed((w2_rsci_qa_d_mxwt[35:18]));
  assign MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_1_nl
      = nl_MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_1_nl[27:0];
  assign MultLoop_mux1h_66_nl = MUX1HOT_v_18_3_2((readslicef_28_18_10((MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_1_nl))),
      z_out_19_27_10, (z_out_18_157_10[17:0]), {and_2670_cse , and_dcpl_1224 , and_dcpl_1228});
  assign nl_z_out_20 = (MultLoop_mux_325_nl) + (MultLoop_mux1h_66_nl);
  assign z_out_20 = nl_z_out_20[17:0];
  assign MultLoop_mux1h_67_nl = MUX1HOT_v_18_3_2((z_out_17[27:10]), (z_out_18_157_10[17:0]),
      z_out_19_27_10, {and_2670_cse , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_21 = ({reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_reg
      , reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_1_reg})
      + (MultLoop_mux1h_67_nl);
  assign z_out_21 = nl_z_out_21[17:0];
  assign nl_ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_sdt
      = conv_s2u_18_19({ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_2_cse
      , ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_19_cse
      , ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_10_cse
      , ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_10_cse})
      + conv_s2u_16_19({ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_2_cse
      , ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_19_cse});
  assign ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_sdt
      = nl_ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_sdt[18:0];
  assign operator_18_8_true_AC_TRN_AC_WRAP_1_mux1h_5_nl = MUX1HOT_s_1_74_2((~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg[2])),
      (~ (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_0_sva_1[17])),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_63_1_ftd),
      (~ (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_63_sva[17])),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_1_ftd),
      (~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_61_1_sva_2[17])),
      (~ (reg_MultLoop_1_mux_64_itm_1_reg[5])), (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_1_ftd),
      (~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_6_1_sva_2[17])),
      (~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_59_1_sva_2[17])),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_1_ftd),
      (~ (reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_reg[5])),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd),
      (~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2[17])),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_1_ftd[2])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd[2])),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_1_ftd),
      (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_1_ftd),
      (~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_58_1_sva_2[17])),
      (~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_60_1_sva_2[17])),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg[2]),
      (reg_MultLoop_1_mux_64_itm_1_reg[5]), (reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_reg[5]),
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_1_ftd,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_1_ftd,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_1_ftd,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd,
      reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd,
      (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2[17]),
      {and_dcpl_1283 , and_dcpl_1289 , and_dcpl_1293 , and_dcpl_1297 , and_dcpl_1301
      , and_dcpl_1302 , and_dcpl_1304 , and_dcpl_1309 , and_dcpl_1313 , and_dcpl_1316
      , and_dcpl_1319 , and_dcpl_1323 , and_dcpl_1325 , and_dcpl_1328 , and_dcpl_1331
      , and_dcpl_1334 , and_dcpl_1339 , and_dcpl_1342 , and_dcpl_1346 , and_dcpl_1350
      , and_dcpl_1353 , and_dcpl_1356 , and_dcpl_1359 , and_dcpl_1362 , and_dcpl_1364
      , and_dcpl_1366 , and_dcpl_1369 , and_dcpl_1371 , and_dcpl_1374 , and_dcpl_1376
      , and_dcpl_1378 , and_dcpl_1380 , and_dcpl_1381 , and_dcpl_1385 , and_dcpl_1387
      , and_dcpl_1389 , and_dcpl_1391 , and_dcpl_1393 , and_dcpl_1395 , and_dcpl_1398
      , and_dcpl_1401 , and_dcpl_1404 , and_dcpl_1406 , and_dcpl_1408 , and_dcpl_1410
      , and_dcpl_1412 , and_dcpl_1413 , and_dcpl_1417 , and_dcpl_1419 , and_dcpl_1421
      , and_dcpl_1423 , and_dcpl_1425 , and_dcpl_1427 , and_dcpl_1429 , and_dcpl_1432
      , and_dcpl_1434 , and_dcpl_1436 , and_dcpl_1438 , and_dcpl_1440 , and_dcpl_1442
      , and_dcpl_1444 , and_dcpl_1445 , and_dcpl_1449 , and_dcpl_1451 , and_1173_cse
      , and_1175_cse , and_1178_cse , and_1180_cse , and_1183_cse , and_1185_cse
      , and_1187_cse , and_1189_cse , and_dcpl_1474 , and_dcpl_1476});
  assign operator_18_8_true_AC_TRN_AC_WRAP_1_mux1h_6_nl = MUX1HOT_v_4_74_2((signext_4_1(~
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg[2]))),
      (signext_4_1(~ (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_0_sva_1[17]))),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_63_1_ftd)),
      (signext_4_1(~ (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_63_sva[17]))),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_1_ftd)),
      (signext_4_1(~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_61_1_sva_2[17]))),
      (signext_4_1(~ (reg_MultLoop_1_mux_64_itm_1_reg[5]))), (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_1_ftd)),
      (signext_4_1(~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_6_1_sva_2[17]))),
      (signext_4_1(~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_59_1_sva_2[17]))),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_1_ftd)),
      (signext_4_1(~ (reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_reg[5]))),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd)),
      (signext_4_1(~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2[17]))),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd)),
      (signext_4_1(~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_1_ftd[2]))),
      (signext_4_1(~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd[2]))),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_1_ftd)),
      (signext_4_1(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_1_ftd)),
      (signext_4_1(~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_58_1_sva_2[17]))),
      (signext_4_1(~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_60_1_sva_2[17]))),
      (nnet_softmax_layer6_t_result_t_softmax_config7_for_1_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_psp_sva_1[14:11]),
      ({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_2_reg
      , reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_4_reg}),
      ({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_1_reg
      , (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_2_reg[11])}),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_14_0[14:11]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_14_0[14:11]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_14_0[14:11]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_14_0[14:11]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_14_0[14:11]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_14_0[14:11]),
      ({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_2_reg
      , (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg[11])}),
      {and_dcpl_1283 , and_dcpl_1289 , and_dcpl_1293 , and_dcpl_1297 , and_dcpl_1301
      , and_dcpl_1302 , and_dcpl_1304 , and_dcpl_1309 , and_dcpl_1313 , and_dcpl_1316
      , and_dcpl_1319 , and_dcpl_1323 , and_dcpl_1325 , and_dcpl_1328 , and_dcpl_1331
      , and_dcpl_1334 , and_dcpl_1339 , and_dcpl_1342 , and_dcpl_1346 , and_dcpl_1350
      , and_dcpl_1353 , and_dcpl_1356 , and_dcpl_1359 , and_dcpl_1362 , and_dcpl_1364
      , and_dcpl_1366 , and_dcpl_1369 , and_dcpl_1371 , and_dcpl_1374 , and_dcpl_1376
      , and_dcpl_1378 , and_dcpl_1380 , and_dcpl_1381 , and_dcpl_1385 , and_dcpl_1387
      , and_dcpl_1389 , and_dcpl_1391 , and_dcpl_1393 , and_dcpl_1395 , and_dcpl_1398
      , and_dcpl_1401 , and_dcpl_1404 , and_dcpl_1406 , and_dcpl_1408 , and_dcpl_1410
      , and_dcpl_1412 , and_dcpl_1413 , and_dcpl_1417 , and_dcpl_1419 , and_dcpl_1421
      , and_dcpl_1423 , and_dcpl_1425 , and_dcpl_1427 , and_dcpl_1429 , and_dcpl_1432
      , and_dcpl_1434 , and_dcpl_1436 , and_dcpl_1438 , and_dcpl_1440 , and_dcpl_1442
      , and_dcpl_1444 , and_dcpl_1445 , and_dcpl_1449 , and_dcpl_1451 , and_1173_cse
      , and_1175_cse , and_1178_cse , and_1180_cse , and_1183_cse , and_1185_cse
      , and_1187_cse , and_1189_cse , and_dcpl_1474 , and_dcpl_1476});
  assign operator_18_8_true_AC_TRN_AC_WRAP_1_mux1h_7_nl = MUX1HOT_v_13_74_2(({(~
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_reg[1:0]))
      , (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_1_reg)
      , (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_2_reg[11:4]))}),
      (~ (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_0_sva_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_63_1_ftd_1[16:4])),
      (~ (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_63_sva[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_1_ftd_1[16:4])),
      (~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_61_1_sva_2[16:4])),
      ({(~ (reg_MultLoop_1_mux_64_itm_1_reg[4:0])) , (~ (reg_MultLoop_1_mux_64_itm_1_1_reg[11:4]))}),
      ({(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_16_15)
      , (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_14_0[14:4]))}),
      ({(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_16_15)
      , (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_14_0[14:4]))}),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_1_ftd_1[16:4])),
      (~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_6_1_sva_2[16:4])),
      (~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_59_1_sva_2[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_1_ftd_1[16:4])),
      ({(~ (reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_reg[4:0]))
      , (~ (reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_1_reg[11:4]))}),
      ({(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_2_reg)
      , (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_4_reg)
      , (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd_2[9:4]))}),
      ({(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_2_reg)
      , (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_3_reg[11:4]))}),
      ({(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_2_reg)
      , (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_3_reg[11:4]))}),
      ({(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_2_reg)
      , (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_3_reg[11:4]))}),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd_1[16:4])),
      (~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2[16:4])),
      ({(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_16_15)
      , (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_14_0[14:4]))}),
      ({(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_16_15)
      , (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_14_0[14:4]))}),
      ({(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_16_15)
      , (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_14_0[14:4]))}),
      ({(~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_16_15)
      , (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_14_0[14:4]))}),
      ({(~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_1_ftd[1:0]))
      , (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_2_reg)
      , (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg[11:4]))}),
      ({(~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd[1:0]))
      , (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_2_reg)
      , (~ reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_4_reg)
      , (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2[10:4]))}),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_1_ftd_1[16:4])),
      (~ (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_1_ftd_1[16:4])),
      (~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_58_1_sva_2[16:4])),
      (~ (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_60_1_sva_2[16:4])),
      ({(nnet_softmax_layer6_t_result_t_softmax_config7_for_1_nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_psp_sva_1[10:0])
      , nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_1_sva_1 , nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_1_sva_1}),
      ({reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2
      , MultLoop_2_and_5_itm_1 , MultLoop_2_and_5_itm_1}), ({(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_2_reg[10:0])
      , MultLoop_2_and_6_itm_1 , MultLoop_2_and_6_itm_1}), ({(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_14_0[10:0])
      , MultLoop_2_and_7_itm_1 , MultLoop_2_and_7_itm_1}), ({(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_14_0[10:0])
      , nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_5_sva , nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_5_sva}),
      ({(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_14_0[10:0])
      , nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_6_sva , nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_6_sva}),
      ({(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_14_0[10:0])
      , nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_7_sva , nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_7_sva}),
      ({(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_14_0[10:0])
      , nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_8_sva , nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_8_sva}),
      ({(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_14_0[10:0])
      , nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_9_sva , nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_9_sva}),
      ({(reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg[10:0])
      , nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_sva , nnet_softmax_layer6_t_result_t_softmax_config7_for_nor_ovfl_sva}),
      {and_dcpl_1283 , and_dcpl_1289 , and_dcpl_1293 , and_dcpl_1297 , and_dcpl_1301
      , and_dcpl_1302 , and_dcpl_1304 , and_dcpl_1309 , and_dcpl_1313 , and_dcpl_1316
      , and_dcpl_1319 , and_dcpl_1323 , and_dcpl_1325 , and_dcpl_1328 , and_dcpl_1331
      , and_dcpl_1334 , and_dcpl_1339 , and_dcpl_1342 , and_dcpl_1346 , and_dcpl_1350
      , and_dcpl_1353 , and_dcpl_1356 , and_dcpl_1359 , and_dcpl_1362 , and_dcpl_1364
      , and_dcpl_1366 , and_dcpl_1369 , and_dcpl_1371 , and_dcpl_1374 , and_dcpl_1376
      , and_dcpl_1378 , and_dcpl_1380 , and_dcpl_1381 , and_dcpl_1385 , and_dcpl_1387
      , and_dcpl_1389 , and_dcpl_1391 , and_dcpl_1393 , and_dcpl_1395 , and_dcpl_1398
      , and_dcpl_1401 , and_dcpl_1404 , and_dcpl_1406 , and_dcpl_1408 , and_dcpl_1410
      , and_dcpl_1412 , and_dcpl_1413 , and_dcpl_1417 , and_dcpl_1419 , and_dcpl_1421
      , and_dcpl_1423 , and_dcpl_1425 , and_dcpl_1427 , and_dcpl_1429 , and_dcpl_1432
      , and_dcpl_1434 , and_dcpl_1436 , and_dcpl_1438 , and_dcpl_1440 , and_dcpl_1442
      , and_dcpl_1444 , and_dcpl_1445 , and_dcpl_1449 , and_dcpl_1451 , and_1173_cse
      , and_1175_cse , and_1178_cse , and_1180_cse , and_1183_cse , and_1185_cse
      , and_1187_cse , and_1189_cse , and_dcpl_1474 , and_dcpl_1476});
  assign operator_18_8_true_AC_TRN_AC_WRAP_1_mux1h_8_nl = MUX1HOT_v_4_64_2((reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_0_1_2_reg[3:0]),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_0_sva_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_63_1_ftd_1[3:0]),
      (nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_acc_63_sva[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_62_1_1_ftd_1[3:0]),
      (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_61_1_sva_2[3:0]),
      (reg_MultLoop_1_mux_64_itm_1_1_reg[3:0]), (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_2_1_1_ftd_1_14_0[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_19_1_1_ftd_1_14_0[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_3_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_29_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_4_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_39_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_5_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_49_1_1_ftd_1[3:0]),
      (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_6_1_sva_2[3:0]),
      (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_59_1_sva_2[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_7_1_1_ftd_1[3:0]),
      (reg_MultLoop_1_2_slc_nnet_dense_large_rf_gt_nin_rem0_layer3_t_layer4_t_config4_MultLoop_1_mux_itm_1_1_reg[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_11_1_1_ftd_2[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_12_1_3_reg[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_13_1_3_reg[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_14_1_3_reg[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_15_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_16_1_1_ftd_1[3:0]),
      (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_17_1_sva_2[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_18_1_1_ftd_1_14_0[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_20_1_1_ftd_1_14_0[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_21_1_1_ftd_1_14_0[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_22_1_1_ftd_1_14_0[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_23_1_3_reg[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_24_1_1_ftd_2[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_25_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_26_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_27_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_28_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_30_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_31_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_32_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_33_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_34_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_35_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_36_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_37_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_38_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_40_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_41_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_42_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_43_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_44_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_45_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_46_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_47_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_48_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_50_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_51_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_52_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_53_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_54_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_55_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_56_1_1_ftd_1[3:0]),
      (reg_nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_57_1_1_ftd_1[3:0]),
      (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_58_1_sva_2[3:0]),
      (nnet_dense_large_rf_gt_nin_rem0_input_t_layer2_t_config2_acc_60_1_sva_2[3:0]),
      {and_dcpl_1283 , and_dcpl_1289 , and_dcpl_1293 , and_dcpl_1297 , and_dcpl_1301
      , and_dcpl_1302 , and_dcpl_1304 , and_dcpl_1309 , and_dcpl_1313 , and_dcpl_1316
      , and_dcpl_1319 , and_dcpl_1323 , and_dcpl_1325 , and_dcpl_1328 , and_dcpl_1331
      , and_dcpl_1334 , and_dcpl_1339 , and_dcpl_1342 , and_dcpl_1346 , and_dcpl_1350
      , and_dcpl_1353 , and_dcpl_1356 , and_dcpl_1359 , and_dcpl_1362 , and_dcpl_1364
      , and_dcpl_1366 , and_dcpl_1369 , and_dcpl_1371 , and_dcpl_1374 , and_dcpl_1376
      , and_dcpl_1378 , and_dcpl_1380 , and_dcpl_1381 , and_dcpl_1385 , and_dcpl_1387
      , and_dcpl_1389 , and_dcpl_1391 , and_dcpl_1393 , and_dcpl_1395 , and_dcpl_1398
      , and_dcpl_1401 , and_dcpl_1404 , and_dcpl_1406 , and_dcpl_1408 , and_dcpl_1410
      , and_dcpl_1412 , and_dcpl_1413 , and_dcpl_1417 , and_dcpl_1419 , and_dcpl_1421
      , and_dcpl_1423 , and_dcpl_1425 , and_dcpl_1427 , and_dcpl_1429 , and_dcpl_1432
      , and_dcpl_1434 , and_dcpl_1436 , and_dcpl_1438 , and_dcpl_1440 , and_dcpl_1442
      , and_dcpl_1444 , and_dcpl_1445 , and_dcpl_1449 , and_dcpl_1451});
  assign operator_18_8_true_AC_TRN_AC_WRAP_1_nor_1_nl = ~(MUX_v_4_2_2((operator_18_8_true_AC_TRN_AC_WRAP_1_mux1h_8_nl),
      4'b1111, operator_18_8_true_AC_TRN_AC_WRAP_1_or_itm));
  assign nl_ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_79_nl
      = conv_s2u_18_19({ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_2_cse
      , ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_19_cse
      , ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_10_cse
      , ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_mux1h_10_cse})
      + conv_s2u_17_19(ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_sdt[18:2]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_79_nl
      = nl_ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_79_nl[18:0];
  assign operator_18_8_true_AC_TRN_AC_WRAP_1_operator_18_8_true_AC_TRN_AC_WRAP_1_operator_18_8_true_AC_TRN_AC_WRAP_1_and_nl
      = MUX_v_19_2_2(19'b0000000000000000000, (ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_79_nl),
      operator_18_8_true_AC_TRN_AC_WRAP_1_or_itm);
  assign operator_18_8_true_AC_TRN_AC_WRAP_1_operator_18_8_true_AC_TRN_AC_WRAP_1_mux_1_nl
      = MUX_v_2_2_2(2'b01, (ac_math_ac_exp_pwl_0_AC_TRN_18_6_true_AC_TRN_AC_SAT_67_47_AC_TRN_AC_WRAP_acc_sdt[1:0]),
      operator_18_8_true_AC_TRN_AC_WRAP_1_or_itm);
  assign nl_operator_18_8_true_AC_TRN_AC_WRAP_1_acc_nl = conv_s2u_22_23({(operator_18_8_true_AC_TRN_AC_WRAP_1_mux1h_5_nl)
      , (operator_18_8_true_AC_TRN_AC_WRAP_1_mux1h_6_nl) , (operator_18_8_true_AC_TRN_AC_WRAP_1_mux1h_7_nl)
      , (operator_18_8_true_AC_TRN_AC_WRAP_1_nor_1_nl)}) + conv_s2u_21_23({(operator_18_8_true_AC_TRN_AC_WRAP_1_operator_18_8_true_AC_TRN_AC_WRAP_1_operator_18_8_true_AC_TRN_AC_WRAP_1_and_nl)
      , (operator_18_8_true_AC_TRN_AC_WRAP_1_operator_18_8_true_AC_TRN_AC_WRAP_1_mux_1_nl)});
  assign operator_18_8_true_AC_TRN_AC_WRAP_1_acc_nl = nl_operator_18_8_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign z_out_23_22_8 = readslicef_23_15_8((operator_18_8_true_AC_TRN_AC_WRAP_1_acc_nl));
  assign SUM_EXP_LOOP_SUM_EXP_LOOP_and_8_nl = (SUM_EXP_LOOP_acc_itm_67_0[67]) & SUM_EXP_LOOP_nor_2_itm;
  assign SUM_EXP_LOOP_mux1h_6_nl = MUX1HOT_v_67_5_2(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_10_18_6_true_AC_TRN_AC_SAT_18_2_AC_TRN_AC_SAT_exp_arr_0_sva,
      CALC_EXP_LOOP_3_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva, CALC_EXP_LOOP_7_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva,
      (SUM_EXP_LOOP_acc_itm_67_0[66:0]), CALC_EXP_LOOP_5_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva,
      {and_dcpl_1483 , and_1282_cse , and_1193_cse , and_1134_cse , and_1286_cse});
  assign SUM_EXP_LOOP_SUM_EXP_LOOP_and_9_nl = (SUM_EXP_LOOP_acc_10_sdt[67]) & SUM_EXP_LOOP_nor_2_itm;
  assign SUM_EXP_LOOP_mux1h_7_nl = MUX1HOT_v_67_5_2(CALC_EXP_LOOP_2_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva,
      CALC_EXP_LOOP_4_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva, CALC_EXP_LOOP_8_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva,
      (SUM_EXP_LOOP_acc_10_sdt[66:0]), CALC_EXP_LOOP_6_operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva,
      {and_dcpl_1483 , and_1282_cse , and_1193_cse , and_1134_cse , and_1286_cse});
  assign nl_z_out_24 = conv_u2u_68_69({(SUM_EXP_LOOP_SUM_EXP_LOOP_and_8_nl) , (SUM_EXP_LOOP_mux1h_6_nl)})
      + conv_u2u_68_69({(SUM_EXP_LOOP_SUM_EXP_LOOP_and_9_nl) , (SUM_EXP_LOOP_mux1h_7_nl)});
  assign z_out_24 = nl_z_out_24[68:0];
  assign mux_1250_nl = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, z_out_12[12:11]);
  assign mux_1249_nl = MUX_v_3_4_2(3'b010, 3'b110, 3'b001, 3'b101, z_out_12[12:11]);
  assign z_out_25 = conv_u2u_19_19(({(mux_1250_nl) , 1'b0 , (mux_1249_nl)}) * (z_out_12[10:1]));

  function automatic [0:0] MUX1HOT_s_1_10_2;
    input [0:0] input_9;
    input [0:0] input_8;
    input [0:0] input_7;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [9:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    result = result | ( input_7 & {1{sel[7]}});
    result = result | ( input_8 & {1{sel[8]}});
    result = result | ( input_9 & {1{sel[9]}});
    MUX1HOT_s_1_10_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_11_2;
    input [0:0] input_10;
    input [0:0] input_9;
    input [0:0] input_8;
    input [0:0] input_7;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [10:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    result = result | ( input_7 & {1{sel[7]}});
    result = result | ( input_8 & {1{sel[8]}});
    result = result | ( input_9 & {1{sel[9]}});
    result = result | ( input_10 & {1{sel[10]}});
    MUX1HOT_s_1_11_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_5_2;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [4:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_74_2;
    input [0:0] input_73;
    input [0:0] input_72;
    input [0:0] input_71;
    input [0:0] input_70;
    input [0:0] input_69;
    input [0:0] input_68;
    input [0:0] input_67;
    input [0:0] input_66;
    input [0:0] input_65;
    input [0:0] input_64;
    input [0:0] input_63;
    input [0:0] input_62;
    input [0:0] input_61;
    input [0:0] input_60;
    input [0:0] input_59;
    input [0:0] input_58;
    input [0:0] input_57;
    input [0:0] input_56;
    input [0:0] input_55;
    input [0:0] input_54;
    input [0:0] input_53;
    input [0:0] input_52;
    input [0:0] input_51;
    input [0:0] input_50;
    input [0:0] input_49;
    input [0:0] input_48;
    input [0:0] input_47;
    input [0:0] input_46;
    input [0:0] input_45;
    input [0:0] input_44;
    input [0:0] input_43;
    input [0:0] input_42;
    input [0:0] input_41;
    input [0:0] input_40;
    input [0:0] input_39;
    input [0:0] input_38;
    input [0:0] input_37;
    input [0:0] input_36;
    input [0:0] input_35;
    input [0:0] input_34;
    input [0:0] input_33;
    input [0:0] input_32;
    input [0:0] input_31;
    input [0:0] input_30;
    input [0:0] input_29;
    input [0:0] input_28;
    input [0:0] input_27;
    input [0:0] input_26;
    input [0:0] input_25;
    input [0:0] input_24;
    input [0:0] input_23;
    input [0:0] input_22;
    input [0:0] input_21;
    input [0:0] input_20;
    input [0:0] input_19;
    input [0:0] input_18;
    input [0:0] input_17;
    input [0:0] input_16;
    input [0:0] input_15;
    input [0:0] input_14;
    input [0:0] input_13;
    input [0:0] input_12;
    input [0:0] input_11;
    input [0:0] input_10;
    input [0:0] input_9;
    input [0:0] input_8;
    input [0:0] input_7;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [73:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    result = result | ( input_7 & {1{sel[7]}});
    result = result | ( input_8 & {1{sel[8]}});
    result = result | ( input_9 & {1{sel[9]}});
    result = result | ( input_10 & {1{sel[10]}});
    result = result | ( input_11 & {1{sel[11]}});
    result = result | ( input_12 & {1{sel[12]}});
    result = result | ( input_13 & {1{sel[13]}});
    result = result | ( input_14 & {1{sel[14]}});
    result = result | ( input_15 & {1{sel[15]}});
    result = result | ( input_16 & {1{sel[16]}});
    result = result | ( input_17 & {1{sel[17]}});
    result = result | ( input_18 & {1{sel[18]}});
    result = result | ( input_19 & {1{sel[19]}});
    result = result | ( input_20 & {1{sel[20]}});
    result = result | ( input_21 & {1{sel[21]}});
    result = result | ( input_22 & {1{sel[22]}});
    result = result | ( input_23 & {1{sel[23]}});
    result = result | ( input_24 & {1{sel[24]}});
    result = result | ( input_25 & {1{sel[25]}});
    result = result | ( input_26 & {1{sel[26]}});
    result = result | ( input_27 & {1{sel[27]}});
    result = result | ( input_28 & {1{sel[28]}});
    result = result | ( input_29 & {1{sel[29]}});
    result = result | ( input_30 & {1{sel[30]}});
    result = result | ( input_31 & {1{sel[31]}});
    result = result | ( input_32 & {1{sel[32]}});
    result = result | ( input_33 & {1{sel[33]}});
    result = result | ( input_34 & {1{sel[34]}});
    result = result | ( input_35 & {1{sel[35]}});
    result = result | ( input_36 & {1{sel[36]}});
    result = result | ( input_37 & {1{sel[37]}});
    result = result | ( input_38 & {1{sel[38]}});
    result = result | ( input_39 & {1{sel[39]}});
    result = result | ( input_40 & {1{sel[40]}});
    result = result | ( input_41 & {1{sel[41]}});
    result = result | ( input_42 & {1{sel[42]}});
    result = result | ( input_43 & {1{sel[43]}});
    result = result | ( input_44 & {1{sel[44]}});
    result = result | ( input_45 & {1{sel[45]}});
    result = result | ( input_46 & {1{sel[46]}});
    result = result | ( input_47 & {1{sel[47]}});
    result = result | ( input_48 & {1{sel[48]}});
    result = result | ( input_49 & {1{sel[49]}});
    result = result | ( input_50 & {1{sel[50]}});
    result = result | ( input_51 & {1{sel[51]}});
    result = result | ( input_52 & {1{sel[52]}});
    result = result | ( input_53 & {1{sel[53]}});
    result = result | ( input_54 & {1{sel[54]}});
    result = result | ( input_55 & {1{sel[55]}});
    result = result | ( input_56 & {1{sel[56]}});
    result = result | ( input_57 & {1{sel[57]}});
    result = result | ( input_58 & {1{sel[58]}});
    result = result | ( input_59 & {1{sel[59]}});
    result = result | ( input_60 & {1{sel[60]}});
    result = result | ( input_61 & {1{sel[61]}});
    result = result | ( input_62 & {1{sel[62]}});
    result = result | ( input_63 & {1{sel[63]}});
    result = result | ( input_64 & {1{sel[64]}});
    result = result | ( input_65 & {1{sel[65]}});
    result = result | ( input_66 & {1{sel[66]}});
    result = result | ( input_67 & {1{sel[67]}});
    result = result | ( input_68 & {1{sel[68]}});
    result = result | ( input_69 & {1{sel[69]}});
    result = result | ( input_70 & {1{sel[70]}});
    result = result | ( input_71 & {1{sel[71]}});
    result = result | ( input_72 & {1{sel[72]}});
    result = result | ( input_73 & {1{sel[73]}});
    MUX1HOT_s_1_74_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_3_2;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [2:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    MUX1HOT_v_10_3_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_9_2;
    input [9:0] input_8;
    input [9:0] input_7;
    input [9:0] input_6;
    input [9:0] input_5;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [8:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    result = result | ( input_3 & {10{sel[3]}});
    result = result | ( input_4 & {10{sel[4]}});
    result = result | ( input_5 & {10{sel[5]}});
    result = result | ( input_6 & {10{sel[6]}});
    result = result | ( input_7 & {10{sel[7]}});
    result = result | ( input_8 & {10{sel[8]}});
    MUX1HOT_v_10_9_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_8_2;
    input [10:0] input_7;
    input [10:0] input_6;
    input [10:0] input_5;
    input [10:0] input_4;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [7:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | ( input_1 & {11{sel[1]}});
    result = result | ( input_2 & {11{sel[2]}});
    result = result | ( input_3 & {11{sel[3]}});
    result = result | ( input_4 & {11{sel[4]}});
    result = result | ( input_5 & {11{sel[5]}});
    result = result | ( input_6 & {11{sel[6]}});
    result = result | ( input_7 & {11{sel[7]}});
    MUX1HOT_v_11_8_2 = result;
  end
  endfunction


  function automatic [11:0] MUX1HOT_v_12_4_2;
    input [11:0] input_3;
    input [11:0] input_2;
    input [11:0] input_1;
    input [11:0] input_0;
    input [3:0] sel;
    reg [11:0] result;
  begin
    result = input_0 & {12{sel[0]}};
    result = result | ( input_1 & {12{sel[1]}});
    result = result | ( input_2 & {12{sel[2]}});
    result = result | ( input_3 & {12{sel[3]}});
    MUX1HOT_v_12_4_2 = result;
  end
  endfunction


  function automatic [12:0] MUX1HOT_v_13_74_2;
    input [12:0] input_73;
    input [12:0] input_72;
    input [12:0] input_71;
    input [12:0] input_70;
    input [12:0] input_69;
    input [12:0] input_68;
    input [12:0] input_67;
    input [12:0] input_66;
    input [12:0] input_65;
    input [12:0] input_64;
    input [12:0] input_63;
    input [12:0] input_62;
    input [12:0] input_61;
    input [12:0] input_60;
    input [12:0] input_59;
    input [12:0] input_58;
    input [12:0] input_57;
    input [12:0] input_56;
    input [12:0] input_55;
    input [12:0] input_54;
    input [12:0] input_53;
    input [12:0] input_52;
    input [12:0] input_51;
    input [12:0] input_50;
    input [12:0] input_49;
    input [12:0] input_48;
    input [12:0] input_47;
    input [12:0] input_46;
    input [12:0] input_45;
    input [12:0] input_44;
    input [12:0] input_43;
    input [12:0] input_42;
    input [12:0] input_41;
    input [12:0] input_40;
    input [12:0] input_39;
    input [12:0] input_38;
    input [12:0] input_37;
    input [12:0] input_36;
    input [12:0] input_35;
    input [12:0] input_34;
    input [12:0] input_33;
    input [12:0] input_32;
    input [12:0] input_31;
    input [12:0] input_30;
    input [12:0] input_29;
    input [12:0] input_28;
    input [12:0] input_27;
    input [12:0] input_26;
    input [12:0] input_25;
    input [12:0] input_24;
    input [12:0] input_23;
    input [12:0] input_22;
    input [12:0] input_21;
    input [12:0] input_20;
    input [12:0] input_19;
    input [12:0] input_18;
    input [12:0] input_17;
    input [12:0] input_16;
    input [12:0] input_15;
    input [12:0] input_14;
    input [12:0] input_13;
    input [12:0] input_12;
    input [12:0] input_11;
    input [12:0] input_10;
    input [12:0] input_9;
    input [12:0] input_8;
    input [12:0] input_7;
    input [12:0] input_6;
    input [12:0] input_5;
    input [12:0] input_4;
    input [12:0] input_3;
    input [12:0] input_2;
    input [12:0] input_1;
    input [12:0] input_0;
    input [73:0] sel;
    reg [12:0] result;
  begin
    result = input_0 & {13{sel[0]}};
    result = result | ( input_1 & {13{sel[1]}});
    result = result | ( input_2 & {13{sel[2]}});
    result = result | ( input_3 & {13{sel[3]}});
    result = result | ( input_4 & {13{sel[4]}});
    result = result | ( input_5 & {13{sel[5]}});
    result = result | ( input_6 & {13{sel[6]}});
    result = result | ( input_7 & {13{sel[7]}});
    result = result | ( input_8 & {13{sel[8]}});
    result = result | ( input_9 & {13{sel[9]}});
    result = result | ( input_10 & {13{sel[10]}});
    result = result | ( input_11 & {13{sel[11]}});
    result = result | ( input_12 & {13{sel[12]}});
    result = result | ( input_13 & {13{sel[13]}});
    result = result | ( input_14 & {13{sel[14]}});
    result = result | ( input_15 & {13{sel[15]}});
    result = result | ( input_16 & {13{sel[16]}});
    result = result | ( input_17 & {13{sel[17]}});
    result = result | ( input_18 & {13{sel[18]}});
    result = result | ( input_19 & {13{sel[19]}});
    result = result | ( input_20 & {13{sel[20]}});
    result = result | ( input_21 & {13{sel[21]}});
    result = result | ( input_22 & {13{sel[22]}});
    result = result | ( input_23 & {13{sel[23]}});
    result = result | ( input_24 & {13{sel[24]}});
    result = result | ( input_25 & {13{sel[25]}});
    result = result | ( input_26 & {13{sel[26]}});
    result = result | ( input_27 & {13{sel[27]}});
    result = result | ( input_28 & {13{sel[28]}});
    result = result | ( input_29 & {13{sel[29]}});
    result = result | ( input_30 & {13{sel[30]}});
    result = result | ( input_31 & {13{sel[31]}});
    result = result | ( input_32 & {13{sel[32]}});
    result = result | ( input_33 & {13{sel[33]}});
    result = result | ( input_34 & {13{sel[34]}});
    result = result | ( input_35 & {13{sel[35]}});
    result = result | ( input_36 & {13{sel[36]}});
    result = result | ( input_37 & {13{sel[37]}});
    result = result | ( input_38 & {13{sel[38]}});
    result = result | ( input_39 & {13{sel[39]}});
    result = result | ( input_40 & {13{sel[40]}});
    result = result | ( input_41 & {13{sel[41]}});
    result = result | ( input_42 & {13{sel[42]}});
    result = result | ( input_43 & {13{sel[43]}});
    result = result | ( input_44 & {13{sel[44]}});
    result = result | ( input_45 & {13{sel[45]}});
    result = result | ( input_46 & {13{sel[46]}});
    result = result | ( input_47 & {13{sel[47]}});
    result = result | ( input_48 & {13{sel[48]}});
    result = result | ( input_49 & {13{sel[49]}});
    result = result | ( input_50 & {13{sel[50]}});
    result = result | ( input_51 & {13{sel[51]}});
    result = result | ( input_52 & {13{sel[52]}});
    result = result | ( input_53 & {13{sel[53]}});
    result = result | ( input_54 & {13{sel[54]}});
    result = result | ( input_55 & {13{sel[55]}});
    result = result | ( input_56 & {13{sel[56]}});
    result = result | ( input_57 & {13{sel[57]}});
    result = result | ( input_58 & {13{sel[58]}});
    result = result | ( input_59 & {13{sel[59]}});
    result = result | ( input_60 & {13{sel[60]}});
    result = result | ( input_61 & {13{sel[61]}});
    result = result | ( input_62 & {13{sel[62]}});
    result = result | ( input_63 & {13{sel[63]}});
    result = result | ( input_64 & {13{sel[64]}});
    result = result | ( input_65 & {13{sel[65]}});
    result = result | ( input_66 & {13{sel[66]}});
    result = result | ( input_67 & {13{sel[67]}});
    result = result | ( input_68 & {13{sel[68]}});
    result = result | ( input_69 & {13{sel[69]}});
    result = result | ( input_70 & {13{sel[70]}});
    result = result | ( input_71 & {13{sel[71]}});
    result = result | ( input_72 & {13{sel[72]}});
    result = result | ( input_73 & {13{sel[73]}});
    MUX1HOT_v_13_74_2 = result;
  end
  endfunction


  function automatic [14:0] MUX1HOT_v_15_10_2;
    input [14:0] input_9;
    input [14:0] input_8;
    input [14:0] input_7;
    input [14:0] input_6;
    input [14:0] input_5;
    input [14:0] input_4;
    input [14:0] input_3;
    input [14:0] input_2;
    input [14:0] input_1;
    input [14:0] input_0;
    input [9:0] sel;
    reg [14:0] result;
  begin
    result = input_0 & {15{sel[0]}};
    result = result | ( input_1 & {15{sel[1]}});
    result = result | ( input_2 & {15{sel[2]}});
    result = result | ( input_3 & {15{sel[3]}});
    result = result | ( input_4 & {15{sel[4]}});
    result = result | ( input_5 & {15{sel[5]}});
    result = result | ( input_6 & {15{sel[6]}});
    result = result | ( input_7 & {15{sel[7]}});
    result = result | ( input_8 & {15{sel[8]}});
    result = result | ( input_9 & {15{sel[9]}});
    MUX1HOT_v_15_10_2 = result;
  end
  endfunction


  function automatic [14:0] MUX1HOT_v_15_11_2;
    input [14:0] input_10;
    input [14:0] input_9;
    input [14:0] input_8;
    input [14:0] input_7;
    input [14:0] input_6;
    input [14:0] input_5;
    input [14:0] input_4;
    input [14:0] input_3;
    input [14:0] input_2;
    input [14:0] input_1;
    input [14:0] input_0;
    input [10:0] sel;
    reg [14:0] result;
  begin
    result = input_0 & {15{sel[0]}};
    result = result | ( input_1 & {15{sel[1]}});
    result = result | ( input_2 & {15{sel[2]}});
    result = result | ( input_3 & {15{sel[3]}});
    result = result | ( input_4 & {15{sel[4]}});
    result = result | ( input_5 & {15{sel[5]}});
    result = result | ( input_6 & {15{sel[6]}});
    result = result | ( input_7 & {15{sel[7]}});
    result = result | ( input_8 & {15{sel[8]}});
    result = result | ( input_9 & {15{sel[9]}});
    result = result | ( input_10 & {15{sel[10]}});
    MUX1HOT_v_15_11_2 = result;
  end
  endfunction


  function automatic [14:0] MUX1HOT_v_15_7_2;
    input [14:0] input_6;
    input [14:0] input_5;
    input [14:0] input_4;
    input [14:0] input_3;
    input [14:0] input_2;
    input [14:0] input_1;
    input [14:0] input_0;
    input [6:0] sel;
    reg [14:0] result;
  begin
    result = input_0 & {15{sel[0]}};
    result = result | ( input_1 & {15{sel[1]}});
    result = result | ( input_2 & {15{sel[2]}});
    result = result | ( input_3 & {15{sel[3]}});
    result = result | ( input_4 & {15{sel[4]}});
    result = result | ( input_5 & {15{sel[5]}});
    result = result | ( input_6 & {15{sel[6]}});
    MUX1HOT_v_15_7_2 = result;
  end
  endfunction


  function automatic [16:0] MUX1HOT_v_17_3_2;
    input [16:0] input_2;
    input [16:0] input_1;
    input [16:0] input_0;
    input [2:0] sel;
    reg [16:0] result;
  begin
    result = input_0 & {17{sel[0]}};
    result = result | ( input_1 & {17{sel[1]}});
    result = result | ( input_2 & {17{sel[2]}});
    MUX1HOT_v_17_3_2 = result;
  end
  endfunction


  function automatic [16:0] MUX1HOT_v_17_6_2;
    input [16:0] input_5;
    input [16:0] input_4;
    input [16:0] input_3;
    input [16:0] input_2;
    input [16:0] input_1;
    input [16:0] input_0;
    input [5:0] sel;
    reg [16:0] result;
  begin
    result = input_0 & {17{sel[0]}};
    result = result | ( input_1 & {17{sel[1]}});
    result = result | ( input_2 & {17{sel[2]}});
    result = result | ( input_3 & {17{sel[3]}});
    result = result | ( input_4 & {17{sel[4]}});
    result = result | ( input_5 & {17{sel[5]}});
    MUX1HOT_v_17_6_2 = result;
  end
  endfunction


  function automatic [16:0] MUX1HOT_v_17_7_2;
    input [16:0] input_6;
    input [16:0] input_5;
    input [16:0] input_4;
    input [16:0] input_3;
    input [16:0] input_2;
    input [16:0] input_1;
    input [16:0] input_0;
    input [6:0] sel;
    reg [16:0] result;
  begin
    result = input_0 & {17{sel[0]}};
    result = result | ( input_1 & {17{sel[1]}});
    result = result | ( input_2 & {17{sel[2]}});
    result = result | ( input_3 & {17{sel[3]}});
    result = result | ( input_4 & {17{sel[4]}});
    result = result | ( input_5 & {17{sel[5]}});
    result = result | ( input_6 & {17{sel[6]}});
    MUX1HOT_v_17_7_2 = result;
  end
  endfunction


  function automatic [16:0] MUX1HOT_v_17_8_2;
    input [16:0] input_7;
    input [16:0] input_6;
    input [16:0] input_5;
    input [16:0] input_4;
    input [16:0] input_3;
    input [16:0] input_2;
    input [16:0] input_1;
    input [16:0] input_0;
    input [7:0] sel;
    reg [16:0] result;
  begin
    result = input_0 & {17{sel[0]}};
    result = result | ( input_1 & {17{sel[1]}});
    result = result | ( input_2 & {17{sel[2]}});
    result = result | ( input_3 & {17{sel[3]}});
    result = result | ( input_4 & {17{sel[4]}});
    result = result | ( input_5 & {17{sel[5]}});
    result = result | ( input_6 & {17{sel[6]}});
    result = result | ( input_7 & {17{sel[7]}});
    MUX1HOT_v_17_8_2 = result;
  end
  endfunction


  function automatic [17:0] MUX1HOT_v_18_12_2;
    input [17:0] input_11;
    input [17:0] input_10;
    input [17:0] input_9;
    input [17:0] input_8;
    input [17:0] input_7;
    input [17:0] input_6;
    input [17:0] input_5;
    input [17:0] input_4;
    input [17:0] input_3;
    input [17:0] input_2;
    input [17:0] input_1;
    input [17:0] input_0;
    input [11:0] sel;
    reg [17:0] result;
  begin
    result = input_0 & {18{sel[0]}};
    result = result | ( input_1 & {18{sel[1]}});
    result = result | ( input_2 & {18{sel[2]}});
    result = result | ( input_3 & {18{sel[3]}});
    result = result | ( input_4 & {18{sel[4]}});
    result = result | ( input_5 & {18{sel[5]}});
    result = result | ( input_6 & {18{sel[6]}});
    result = result | ( input_7 & {18{sel[7]}});
    result = result | ( input_8 & {18{sel[8]}});
    result = result | ( input_9 & {18{sel[9]}});
    result = result | ( input_10 & {18{sel[10]}});
    result = result | ( input_11 & {18{sel[11]}});
    MUX1HOT_v_18_12_2 = result;
  end
  endfunction


  function automatic [17:0] MUX1HOT_v_18_13_2;
    input [17:0] input_12;
    input [17:0] input_11;
    input [17:0] input_10;
    input [17:0] input_9;
    input [17:0] input_8;
    input [17:0] input_7;
    input [17:0] input_6;
    input [17:0] input_5;
    input [17:0] input_4;
    input [17:0] input_3;
    input [17:0] input_2;
    input [17:0] input_1;
    input [17:0] input_0;
    input [12:0] sel;
    reg [17:0] result;
  begin
    result = input_0 & {18{sel[0]}};
    result = result | ( input_1 & {18{sel[1]}});
    result = result | ( input_2 & {18{sel[2]}});
    result = result | ( input_3 & {18{sel[3]}});
    result = result | ( input_4 & {18{sel[4]}});
    result = result | ( input_5 & {18{sel[5]}});
    result = result | ( input_6 & {18{sel[6]}});
    result = result | ( input_7 & {18{sel[7]}});
    result = result | ( input_8 & {18{sel[8]}});
    result = result | ( input_9 & {18{sel[9]}});
    result = result | ( input_10 & {18{sel[10]}});
    result = result | ( input_11 & {18{sel[11]}});
    result = result | ( input_12 & {18{sel[12]}});
    MUX1HOT_v_18_13_2 = result;
  end
  endfunction


  function automatic [17:0] MUX1HOT_v_18_3_2;
    input [17:0] input_2;
    input [17:0] input_1;
    input [17:0] input_0;
    input [2:0] sel;
    reg [17:0] result;
  begin
    result = input_0 & {18{sel[0]}};
    result = result | ( input_1 & {18{sel[1]}});
    result = result | ( input_2 & {18{sel[2]}});
    MUX1HOT_v_18_3_2 = result;
  end
  endfunction


  function automatic [17:0] MUX1HOT_v_18_4_2;
    input [17:0] input_3;
    input [17:0] input_2;
    input [17:0] input_1;
    input [17:0] input_0;
    input [3:0] sel;
    reg [17:0] result;
  begin
    result = input_0 & {18{sel[0]}};
    result = result | ( input_1 & {18{sel[1]}});
    result = result | ( input_2 & {18{sel[2]}});
    result = result | ( input_3 & {18{sel[3]}});
    MUX1HOT_v_18_4_2 = result;
  end
  endfunction


  function automatic [17:0] MUX1HOT_v_18_5_2;
    input [17:0] input_4;
    input [17:0] input_3;
    input [17:0] input_2;
    input [17:0] input_1;
    input [17:0] input_0;
    input [4:0] sel;
    reg [17:0] result;
  begin
    result = input_0 & {18{sel[0]}};
    result = result | ( input_1 & {18{sel[1]}});
    result = result | ( input_2 & {18{sel[2]}});
    result = result | ( input_3 & {18{sel[3]}});
    result = result | ( input_4 & {18{sel[4]}});
    MUX1HOT_v_18_5_2 = result;
  end
  endfunction


  function automatic [17:0] MUX1HOT_v_18_7_2;
    input [17:0] input_6;
    input [17:0] input_5;
    input [17:0] input_4;
    input [17:0] input_3;
    input [17:0] input_2;
    input [17:0] input_1;
    input [17:0] input_0;
    input [6:0] sel;
    reg [17:0] result;
  begin
    result = input_0 & {18{sel[0]}};
    result = result | ( input_1 & {18{sel[1]}});
    result = result | ( input_2 & {18{sel[2]}});
    result = result | ( input_3 & {18{sel[3]}});
    result = result | ( input_4 & {18{sel[4]}});
    result = result | ( input_5 & {18{sel[5]}});
    result = result | ( input_6 & {18{sel[6]}});
    MUX1HOT_v_18_7_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    result = result | ( input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_5_2;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [4:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    result = result | ( input_3 & {3{sel[3]}});
    result = result | ( input_4 & {3{sel[4]}});
    MUX1HOT_v_3_5_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_64_2;
    input [3:0] input_63;
    input [3:0] input_62;
    input [3:0] input_61;
    input [3:0] input_60;
    input [3:0] input_59;
    input [3:0] input_58;
    input [3:0] input_57;
    input [3:0] input_56;
    input [3:0] input_55;
    input [3:0] input_54;
    input [3:0] input_53;
    input [3:0] input_52;
    input [3:0] input_51;
    input [3:0] input_50;
    input [3:0] input_49;
    input [3:0] input_48;
    input [3:0] input_47;
    input [3:0] input_46;
    input [3:0] input_45;
    input [3:0] input_44;
    input [3:0] input_43;
    input [3:0] input_42;
    input [3:0] input_41;
    input [3:0] input_40;
    input [3:0] input_39;
    input [3:0] input_38;
    input [3:0] input_37;
    input [3:0] input_36;
    input [3:0] input_35;
    input [3:0] input_34;
    input [3:0] input_33;
    input [3:0] input_32;
    input [3:0] input_31;
    input [3:0] input_30;
    input [3:0] input_29;
    input [3:0] input_28;
    input [3:0] input_27;
    input [3:0] input_26;
    input [3:0] input_25;
    input [3:0] input_24;
    input [3:0] input_23;
    input [3:0] input_22;
    input [3:0] input_21;
    input [3:0] input_20;
    input [3:0] input_19;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [63:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    result = result | ( input_4 & {4{sel[4]}});
    result = result | ( input_5 & {4{sel[5]}});
    result = result | ( input_6 & {4{sel[6]}});
    result = result | ( input_7 & {4{sel[7]}});
    result = result | ( input_8 & {4{sel[8]}});
    result = result | ( input_9 & {4{sel[9]}});
    result = result | ( input_10 & {4{sel[10]}});
    result = result | ( input_11 & {4{sel[11]}});
    result = result | ( input_12 & {4{sel[12]}});
    result = result | ( input_13 & {4{sel[13]}});
    result = result | ( input_14 & {4{sel[14]}});
    result = result | ( input_15 & {4{sel[15]}});
    result = result | ( input_16 & {4{sel[16]}});
    result = result | ( input_17 & {4{sel[17]}});
    result = result | ( input_18 & {4{sel[18]}});
    result = result | ( input_19 & {4{sel[19]}});
    result = result | ( input_20 & {4{sel[20]}});
    result = result | ( input_21 & {4{sel[21]}});
    result = result | ( input_22 & {4{sel[22]}});
    result = result | ( input_23 & {4{sel[23]}});
    result = result | ( input_24 & {4{sel[24]}});
    result = result | ( input_25 & {4{sel[25]}});
    result = result | ( input_26 & {4{sel[26]}});
    result = result | ( input_27 & {4{sel[27]}});
    result = result | ( input_28 & {4{sel[28]}});
    result = result | ( input_29 & {4{sel[29]}});
    result = result | ( input_30 & {4{sel[30]}});
    result = result | ( input_31 & {4{sel[31]}});
    result = result | ( input_32 & {4{sel[32]}});
    result = result | ( input_33 & {4{sel[33]}});
    result = result | ( input_34 & {4{sel[34]}});
    result = result | ( input_35 & {4{sel[35]}});
    result = result | ( input_36 & {4{sel[36]}});
    result = result | ( input_37 & {4{sel[37]}});
    result = result | ( input_38 & {4{sel[38]}});
    result = result | ( input_39 & {4{sel[39]}});
    result = result | ( input_40 & {4{sel[40]}});
    result = result | ( input_41 & {4{sel[41]}});
    result = result | ( input_42 & {4{sel[42]}});
    result = result | ( input_43 & {4{sel[43]}});
    result = result | ( input_44 & {4{sel[44]}});
    result = result | ( input_45 & {4{sel[45]}});
    result = result | ( input_46 & {4{sel[46]}});
    result = result | ( input_47 & {4{sel[47]}});
    result = result | ( input_48 & {4{sel[48]}});
    result = result | ( input_49 & {4{sel[49]}});
    result = result | ( input_50 & {4{sel[50]}});
    result = result | ( input_51 & {4{sel[51]}});
    result = result | ( input_52 & {4{sel[52]}});
    result = result | ( input_53 & {4{sel[53]}});
    result = result | ( input_54 & {4{sel[54]}});
    result = result | ( input_55 & {4{sel[55]}});
    result = result | ( input_56 & {4{sel[56]}});
    result = result | ( input_57 & {4{sel[57]}});
    result = result | ( input_58 & {4{sel[58]}});
    result = result | ( input_59 & {4{sel[59]}});
    result = result | ( input_60 & {4{sel[60]}});
    result = result | ( input_61 & {4{sel[61]}});
    result = result | ( input_62 & {4{sel[62]}});
    result = result | ( input_63 & {4{sel[63]}});
    MUX1HOT_v_4_64_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_6_2;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [5:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    result = result | ( input_4 & {4{sel[4]}});
    result = result | ( input_5 & {4{sel[5]}});
    MUX1HOT_v_4_6_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_74_2;
    input [3:0] input_73;
    input [3:0] input_72;
    input [3:0] input_71;
    input [3:0] input_70;
    input [3:0] input_69;
    input [3:0] input_68;
    input [3:0] input_67;
    input [3:0] input_66;
    input [3:0] input_65;
    input [3:0] input_64;
    input [3:0] input_63;
    input [3:0] input_62;
    input [3:0] input_61;
    input [3:0] input_60;
    input [3:0] input_59;
    input [3:0] input_58;
    input [3:0] input_57;
    input [3:0] input_56;
    input [3:0] input_55;
    input [3:0] input_54;
    input [3:0] input_53;
    input [3:0] input_52;
    input [3:0] input_51;
    input [3:0] input_50;
    input [3:0] input_49;
    input [3:0] input_48;
    input [3:0] input_47;
    input [3:0] input_46;
    input [3:0] input_45;
    input [3:0] input_44;
    input [3:0] input_43;
    input [3:0] input_42;
    input [3:0] input_41;
    input [3:0] input_40;
    input [3:0] input_39;
    input [3:0] input_38;
    input [3:0] input_37;
    input [3:0] input_36;
    input [3:0] input_35;
    input [3:0] input_34;
    input [3:0] input_33;
    input [3:0] input_32;
    input [3:0] input_31;
    input [3:0] input_30;
    input [3:0] input_29;
    input [3:0] input_28;
    input [3:0] input_27;
    input [3:0] input_26;
    input [3:0] input_25;
    input [3:0] input_24;
    input [3:0] input_23;
    input [3:0] input_22;
    input [3:0] input_21;
    input [3:0] input_20;
    input [3:0] input_19;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [73:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    result = result | ( input_4 & {4{sel[4]}});
    result = result | ( input_5 & {4{sel[5]}});
    result = result | ( input_6 & {4{sel[6]}});
    result = result | ( input_7 & {4{sel[7]}});
    result = result | ( input_8 & {4{sel[8]}});
    result = result | ( input_9 & {4{sel[9]}});
    result = result | ( input_10 & {4{sel[10]}});
    result = result | ( input_11 & {4{sel[11]}});
    result = result | ( input_12 & {4{sel[12]}});
    result = result | ( input_13 & {4{sel[13]}});
    result = result | ( input_14 & {4{sel[14]}});
    result = result | ( input_15 & {4{sel[15]}});
    result = result | ( input_16 & {4{sel[16]}});
    result = result | ( input_17 & {4{sel[17]}});
    result = result | ( input_18 & {4{sel[18]}});
    result = result | ( input_19 & {4{sel[19]}});
    result = result | ( input_20 & {4{sel[20]}});
    result = result | ( input_21 & {4{sel[21]}});
    result = result | ( input_22 & {4{sel[22]}});
    result = result | ( input_23 & {4{sel[23]}});
    result = result | ( input_24 & {4{sel[24]}});
    result = result | ( input_25 & {4{sel[25]}});
    result = result | ( input_26 & {4{sel[26]}});
    result = result | ( input_27 & {4{sel[27]}});
    result = result | ( input_28 & {4{sel[28]}});
    result = result | ( input_29 & {4{sel[29]}});
    result = result | ( input_30 & {4{sel[30]}});
    result = result | ( input_31 & {4{sel[31]}});
    result = result | ( input_32 & {4{sel[32]}});
    result = result | ( input_33 & {4{sel[33]}});
    result = result | ( input_34 & {4{sel[34]}});
    result = result | ( input_35 & {4{sel[35]}});
    result = result | ( input_36 & {4{sel[36]}});
    result = result | ( input_37 & {4{sel[37]}});
    result = result | ( input_38 & {4{sel[38]}});
    result = result | ( input_39 & {4{sel[39]}});
    result = result | ( input_40 & {4{sel[40]}});
    result = result | ( input_41 & {4{sel[41]}});
    result = result | ( input_42 & {4{sel[42]}});
    result = result | ( input_43 & {4{sel[43]}});
    result = result | ( input_44 & {4{sel[44]}});
    result = result | ( input_45 & {4{sel[45]}});
    result = result | ( input_46 & {4{sel[46]}});
    result = result | ( input_47 & {4{sel[47]}});
    result = result | ( input_48 & {4{sel[48]}});
    result = result | ( input_49 & {4{sel[49]}});
    result = result | ( input_50 & {4{sel[50]}});
    result = result | ( input_51 & {4{sel[51]}});
    result = result | ( input_52 & {4{sel[52]}});
    result = result | ( input_53 & {4{sel[53]}});
    result = result | ( input_54 & {4{sel[54]}});
    result = result | ( input_55 & {4{sel[55]}});
    result = result | ( input_56 & {4{sel[56]}});
    result = result | ( input_57 & {4{sel[57]}});
    result = result | ( input_58 & {4{sel[58]}});
    result = result | ( input_59 & {4{sel[59]}});
    result = result | ( input_60 & {4{sel[60]}});
    result = result | ( input_61 & {4{sel[61]}});
    result = result | ( input_62 & {4{sel[62]}});
    result = result | ( input_63 & {4{sel[63]}});
    result = result | ( input_64 & {4{sel[64]}});
    result = result | ( input_65 & {4{sel[65]}});
    result = result | ( input_66 & {4{sel[66]}});
    result = result | ( input_67 & {4{sel[67]}});
    result = result | ( input_68 & {4{sel[68]}});
    result = result | ( input_69 & {4{sel[69]}});
    result = result | ( input_70 & {4{sel[70]}});
    result = result | ( input_71 & {4{sel[71]}});
    result = result | ( input_72 & {4{sel[72]}});
    result = result | ( input_73 & {4{sel[73]}});
    MUX1HOT_v_4_74_2 = result;
  end
  endfunction


  function automatic [66:0] MUX1HOT_v_67_11_2;
    input [66:0] input_10;
    input [66:0] input_9;
    input [66:0] input_8;
    input [66:0] input_7;
    input [66:0] input_6;
    input [66:0] input_5;
    input [66:0] input_4;
    input [66:0] input_3;
    input [66:0] input_2;
    input [66:0] input_1;
    input [66:0] input_0;
    input [10:0] sel;
    reg [66:0] result;
  begin
    result = input_0 & {67{sel[0]}};
    result = result | ( input_1 & {67{sel[1]}});
    result = result | ( input_2 & {67{sel[2]}});
    result = result | ( input_3 & {67{sel[3]}});
    result = result | ( input_4 & {67{sel[4]}});
    result = result | ( input_5 & {67{sel[5]}});
    result = result | ( input_6 & {67{sel[6]}});
    result = result | ( input_7 & {67{sel[7]}});
    result = result | ( input_8 & {67{sel[8]}});
    result = result | ( input_9 & {67{sel[9]}});
    result = result | ( input_10 & {67{sel[10]}});
    MUX1HOT_v_67_11_2 = result;
  end
  endfunction


  function automatic [66:0] MUX1HOT_v_67_5_2;
    input [66:0] input_4;
    input [66:0] input_3;
    input [66:0] input_2;
    input [66:0] input_1;
    input [66:0] input_0;
    input [4:0] sel;
    reg [66:0] result;
  begin
    result = input_0 & {67{sel[0]}};
    result = result | ( input_1 & {67{sel[1]}});
    result = result | ( input_2 & {67{sel[2]}});
    result = result | ( input_3 & {67{sel[3]}});
    result = result | ( input_4 & {67{sel[4]}});
    MUX1HOT_v_67_5_2 = result;
  end
  endfunction


  function automatic [67:0] MUX1HOT_v_68_3_2;
    input [67:0] input_2;
    input [67:0] input_1;
    input [67:0] input_0;
    input [2:0] sel;
    reg [67:0] result;
  begin
    result = input_0 & {68{sel[0]}};
    result = result | ( input_1 & {68{sel[1]}});
    result = result | ( input_2 & {68{sel[2]}});
    MUX1HOT_v_68_3_2 = result;
  end
  endfunction


  function automatic [73:0] MUX1HOT_v_74_3_2;
    input [73:0] input_2;
    input [73:0] input_1;
    input [73:0] input_0;
    input [2:0] sel;
    reg [73:0] result;
  begin
    result = input_0 & {74{sel[0]}};
    result = result | ( input_1 & {74{sel[1]}});
    result = result | ( input_2 & {74{sel[2]}});
    MUX1HOT_v_74_3_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_8_2;
    input [6:0] input_7;
    input [6:0] input_6;
    input [6:0] input_5;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [7:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    result = result | ( input_3 & {7{sel[3]}});
    result = result | ( input_4 & {7{sel[4]}});
    result = result | ( input_5 & {7{sel[5]}});
    result = result | ( input_6 & {7{sel[6]}});
    result = result | ( input_7 & {7{sel[7]}});
    MUX1HOT_v_7_8_2 = result;
  end
  endfunction


  function automatic [8:0] MUX1HOT_v_9_3_2;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [2:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | ( input_1 & {9{sel[1]}});
    result = result | ( input_2 & {9{sel[2]}});
    MUX1HOT_v_9_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_10_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input [11:0] input_2;
    input [11:0] input_3;
    input [11:0] input_4;
    input [11:0] input_5;
    input [11:0] input_6;
    input [11:0] input_7;
    input [11:0] input_8;
    input [11:0] input_9;
    input [3:0] sel;
    reg [11:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      default : begin
        result = input_9;
      end
    endcase
    MUX_v_12_10_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input [0:0] sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [14:0] MUX_v_15_2_2;
    input [14:0] input_0;
    input [14:0] input_1;
    input [0:0] sel;
    reg [14:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_15_2_2 = result;
  end
  endfunction


  function automatic [14:0] MUX_v_15_64_2;
    input [14:0] input_0;
    input [14:0] input_1;
    input [14:0] input_2;
    input [14:0] input_3;
    input [14:0] input_4;
    input [14:0] input_5;
    input [14:0] input_6;
    input [14:0] input_7;
    input [14:0] input_8;
    input [14:0] input_9;
    input [14:0] input_10;
    input [14:0] input_11;
    input [14:0] input_12;
    input [14:0] input_13;
    input [14:0] input_14;
    input [14:0] input_15;
    input [14:0] input_16;
    input [14:0] input_17;
    input [14:0] input_18;
    input [14:0] input_19;
    input [14:0] input_20;
    input [14:0] input_21;
    input [14:0] input_22;
    input [14:0] input_23;
    input [14:0] input_24;
    input [14:0] input_25;
    input [14:0] input_26;
    input [14:0] input_27;
    input [14:0] input_28;
    input [14:0] input_29;
    input [14:0] input_30;
    input [14:0] input_31;
    input [14:0] input_32;
    input [14:0] input_33;
    input [14:0] input_34;
    input [14:0] input_35;
    input [14:0] input_36;
    input [14:0] input_37;
    input [14:0] input_38;
    input [14:0] input_39;
    input [14:0] input_40;
    input [14:0] input_41;
    input [14:0] input_42;
    input [14:0] input_43;
    input [14:0] input_44;
    input [14:0] input_45;
    input [14:0] input_46;
    input [14:0] input_47;
    input [14:0] input_48;
    input [14:0] input_49;
    input [14:0] input_50;
    input [14:0] input_51;
    input [14:0] input_52;
    input [14:0] input_53;
    input [14:0] input_54;
    input [14:0] input_55;
    input [14:0] input_56;
    input [14:0] input_57;
    input [14:0] input_58;
    input [14:0] input_59;
    input [14:0] input_60;
    input [14:0] input_61;
    input [14:0] input_62;
    input [14:0] input_63;
    input [5:0] sel;
    reg [14:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_15_64_2 = result;
  end
  endfunction


  function automatic [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction


  function automatic [17:0] MUX_v_18_10_2;
    input [17:0] input_0;
    input [17:0] input_1;
    input [17:0] input_2;
    input [17:0] input_3;
    input [17:0] input_4;
    input [17:0] input_5;
    input [17:0] input_6;
    input [17:0] input_7;
    input [17:0] input_8;
    input [17:0] input_9;
    input [3:0] sel;
    reg [17:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      default : begin
        result = input_9;
      end
    endcase
    MUX_v_18_10_2 = result;
  end
  endfunction


  function automatic [17:0] MUX_v_18_2_2;
    input [17:0] input_0;
    input [17:0] input_1;
    input [0:0] sel;
    reg [17:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_18_2_2 = result;
  end
  endfunction


  function automatic [17:0] MUX_v_18_32_2;
    input [17:0] input_0;
    input [17:0] input_1;
    input [17:0] input_2;
    input [17:0] input_3;
    input [17:0] input_4;
    input [17:0] input_5;
    input [17:0] input_6;
    input [17:0] input_7;
    input [17:0] input_8;
    input [17:0] input_9;
    input [17:0] input_10;
    input [17:0] input_11;
    input [17:0] input_12;
    input [17:0] input_13;
    input [17:0] input_14;
    input [17:0] input_15;
    input [17:0] input_16;
    input [17:0] input_17;
    input [17:0] input_18;
    input [17:0] input_19;
    input [17:0] input_20;
    input [17:0] input_21;
    input [17:0] input_22;
    input [17:0] input_23;
    input [17:0] input_24;
    input [17:0] input_25;
    input [17:0] input_26;
    input [17:0] input_27;
    input [17:0] input_28;
    input [17:0] input_29;
    input [17:0] input_30;
    input [17:0] input_31;
    input [4:0] sel;
    reg [17:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_v_18_32_2 = result;
  end
  endfunction


  function automatic [17:0] MUX_v_18_64_2;
    input [17:0] input_0;
    input [17:0] input_1;
    input [17:0] input_2;
    input [17:0] input_3;
    input [17:0] input_4;
    input [17:0] input_5;
    input [17:0] input_6;
    input [17:0] input_7;
    input [17:0] input_8;
    input [17:0] input_9;
    input [17:0] input_10;
    input [17:0] input_11;
    input [17:0] input_12;
    input [17:0] input_13;
    input [17:0] input_14;
    input [17:0] input_15;
    input [17:0] input_16;
    input [17:0] input_17;
    input [17:0] input_18;
    input [17:0] input_19;
    input [17:0] input_20;
    input [17:0] input_21;
    input [17:0] input_22;
    input [17:0] input_23;
    input [17:0] input_24;
    input [17:0] input_25;
    input [17:0] input_26;
    input [17:0] input_27;
    input [17:0] input_28;
    input [17:0] input_29;
    input [17:0] input_30;
    input [17:0] input_31;
    input [17:0] input_32;
    input [17:0] input_33;
    input [17:0] input_34;
    input [17:0] input_35;
    input [17:0] input_36;
    input [17:0] input_37;
    input [17:0] input_38;
    input [17:0] input_39;
    input [17:0] input_40;
    input [17:0] input_41;
    input [17:0] input_42;
    input [17:0] input_43;
    input [17:0] input_44;
    input [17:0] input_45;
    input [17:0] input_46;
    input [17:0] input_47;
    input [17:0] input_48;
    input [17:0] input_49;
    input [17:0] input_50;
    input [17:0] input_51;
    input [17:0] input_52;
    input [17:0] input_53;
    input [17:0] input_54;
    input [17:0] input_55;
    input [17:0] input_56;
    input [17:0] input_57;
    input [17:0] input_58;
    input [17:0] input_59;
    input [17:0] input_60;
    input [17:0] input_61;
    input [17:0] input_62;
    input [17:0] input_63;
    input [5:0] sel;
    reg [17:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_18_64_2 = result;
  end
  endfunction


  function automatic [17:0] MUX_v_18_784_2;
    input [17:0] input_0;
    input [17:0] input_1;
    input [17:0] input_2;
    input [17:0] input_3;
    input [17:0] input_4;
    input [17:0] input_5;
    input [17:0] input_6;
    input [17:0] input_7;
    input [17:0] input_8;
    input [17:0] input_9;
    input [17:0] input_10;
    input [17:0] input_11;
    input [17:0] input_12;
    input [17:0] input_13;
    input [17:0] input_14;
    input [17:0] input_15;
    input [17:0] input_16;
    input [17:0] input_17;
    input [17:0] input_18;
    input [17:0] input_19;
    input [17:0] input_20;
    input [17:0] input_21;
    input [17:0] input_22;
    input [17:0] input_23;
    input [17:0] input_24;
    input [17:0] input_25;
    input [17:0] input_26;
    input [17:0] input_27;
    input [17:0] input_28;
    input [17:0] input_29;
    input [17:0] input_30;
    input [17:0] input_31;
    input [17:0] input_32;
    input [17:0] input_33;
    input [17:0] input_34;
    input [17:0] input_35;
    input [17:0] input_36;
    input [17:0] input_37;
    input [17:0] input_38;
    input [17:0] input_39;
    input [17:0] input_40;
    input [17:0] input_41;
    input [17:0] input_42;
    input [17:0] input_43;
    input [17:0] input_44;
    input [17:0] input_45;
    input [17:0] input_46;
    input [17:0] input_47;
    input [17:0] input_48;
    input [17:0] input_49;
    input [17:0] input_50;
    input [17:0] input_51;
    input [17:0] input_52;
    input [17:0] input_53;
    input [17:0] input_54;
    input [17:0] input_55;
    input [17:0] input_56;
    input [17:0] input_57;
    input [17:0] input_58;
    input [17:0] input_59;
    input [17:0] input_60;
    input [17:0] input_61;
    input [17:0] input_62;
    input [17:0] input_63;
    input [17:0] input_64;
    input [17:0] input_65;
    input [17:0] input_66;
    input [17:0] input_67;
    input [17:0] input_68;
    input [17:0] input_69;
    input [17:0] input_70;
    input [17:0] input_71;
    input [17:0] input_72;
    input [17:0] input_73;
    input [17:0] input_74;
    input [17:0] input_75;
    input [17:0] input_76;
    input [17:0] input_77;
    input [17:0] input_78;
    input [17:0] input_79;
    input [17:0] input_80;
    input [17:0] input_81;
    input [17:0] input_82;
    input [17:0] input_83;
    input [17:0] input_84;
    input [17:0] input_85;
    input [17:0] input_86;
    input [17:0] input_87;
    input [17:0] input_88;
    input [17:0] input_89;
    input [17:0] input_90;
    input [17:0] input_91;
    input [17:0] input_92;
    input [17:0] input_93;
    input [17:0] input_94;
    input [17:0] input_95;
    input [17:0] input_96;
    input [17:0] input_97;
    input [17:0] input_98;
    input [17:0] input_99;
    input [17:0] input_100;
    input [17:0] input_101;
    input [17:0] input_102;
    input [17:0] input_103;
    input [17:0] input_104;
    input [17:0] input_105;
    input [17:0] input_106;
    input [17:0] input_107;
    input [17:0] input_108;
    input [17:0] input_109;
    input [17:0] input_110;
    input [17:0] input_111;
    input [17:0] input_112;
    input [17:0] input_113;
    input [17:0] input_114;
    input [17:0] input_115;
    input [17:0] input_116;
    input [17:0] input_117;
    input [17:0] input_118;
    input [17:0] input_119;
    input [17:0] input_120;
    input [17:0] input_121;
    input [17:0] input_122;
    input [17:0] input_123;
    input [17:0] input_124;
    input [17:0] input_125;
    input [17:0] input_126;
    input [17:0] input_127;
    input [17:0] input_128;
    input [17:0] input_129;
    input [17:0] input_130;
    input [17:0] input_131;
    input [17:0] input_132;
    input [17:0] input_133;
    input [17:0] input_134;
    input [17:0] input_135;
    input [17:0] input_136;
    input [17:0] input_137;
    input [17:0] input_138;
    input [17:0] input_139;
    input [17:0] input_140;
    input [17:0] input_141;
    input [17:0] input_142;
    input [17:0] input_143;
    input [17:0] input_144;
    input [17:0] input_145;
    input [17:0] input_146;
    input [17:0] input_147;
    input [17:0] input_148;
    input [17:0] input_149;
    input [17:0] input_150;
    input [17:0] input_151;
    input [17:0] input_152;
    input [17:0] input_153;
    input [17:0] input_154;
    input [17:0] input_155;
    input [17:0] input_156;
    input [17:0] input_157;
    input [17:0] input_158;
    input [17:0] input_159;
    input [17:0] input_160;
    input [17:0] input_161;
    input [17:0] input_162;
    input [17:0] input_163;
    input [17:0] input_164;
    input [17:0] input_165;
    input [17:0] input_166;
    input [17:0] input_167;
    input [17:0] input_168;
    input [17:0] input_169;
    input [17:0] input_170;
    input [17:0] input_171;
    input [17:0] input_172;
    input [17:0] input_173;
    input [17:0] input_174;
    input [17:0] input_175;
    input [17:0] input_176;
    input [17:0] input_177;
    input [17:0] input_178;
    input [17:0] input_179;
    input [17:0] input_180;
    input [17:0] input_181;
    input [17:0] input_182;
    input [17:0] input_183;
    input [17:0] input_184;
    input [17:0] input_185;
    input [17:0] input_186;
    input [17:0] input_187;
    input [17:0] input_188;
    input [17:0] input_189;
    input [17:0] input_190;
    input [17:0] input_191;
    input [17:0] input_192;
    input [17:0] input_193;
    input [17:0] input_194;
    input [17:0] input_195;
    input [17:0] input_196;
    input [17:0] input_197;
    input [17:0] input_198;
    input [17:0] input_199;
    input [17:0] input_200;
    input [17:0] input_201;
    input [17:0] input_202;
    input [17:0] input_203;
    input [17:0] input_204;
    input [17:0] input_205;
    input [17:0] input_206;
    input [17:0] input_207;
    input [17:0] input_208;
    input [17:0] input_209;
    input [17:0] input_210;
    input [17:0] input_211;
    input [17:0] input_212;
    input [17:0] input_213;
    input [17:0] input_214;
    input [17:0] input_215;
    input [17:0] input_216;
    input [17:0] input_217;
    input [17:0] input_218;
    input [17:0] input_219;
    input [17:0] input_220;
    input [17:0] input_221;
    input [17:0] input_222;
    input [17:0] input_223;
    input [17:0] input_224;
    input [17:0] input_225;
    input [17:0] input_226;
    input [17:0] input_227;
    input [17:0] input_228;
    input [17:0] input_229;
    input [17:0] input_230;
    input [17:0] input_231;
    input [17:0] input_232;
    input [17:0] input_233;
    input [17:0] input_234;
    input [17:0] input_235;
    input [17:0] input_236;
    input [17:0] input_237;
    input [17:0] input_238;
    input [17:0] input_239;
    input [17:0] input_240;
    input [17:0] input_241;
    input [17:0] input_242;
    input [17:0] input_243;
    input [17:0] input_244;
    input [17:0] input_245;
    input [17:0] input_246;
    input [17:0] input_247;
    input [17:0] input_248;
    input [17:0] input_249;
    input [17:0] input_250;
    input [17:0] input_251;
    input [17:0] input_252;
    input [17:0] input_253;
    input [17:0] input_254;
    input [17:0] input_255;
    input [17:0] input_256;
    input [17:0] input_257;
    input [17:0] input_258;
    input [17:0] input_259;
    input [17:0] input_260;
    input [17:0] input_261;
    input [17:0] input_262;
    input [17:0] input_263;
    input [17:0] input_264;
    input [17:0] input_265;
    input [17:0] input_266;
    input [17:0] input_267;
    input [17:0] input_268;
    input [17:0] input_269;
    input [17:0] input_270;
    input [17:0] input_271;
    input [17:0] input_272;
    input [17:0] input_273;
    input [17:0] input_274;
    input [17:0] input_275;
    input [17:0] input_276;
    input [17:0] input_277;
    input [17:0] input_278;
    input [17:0] input_279;
    input [17:0] input_280;
    input [17:0] input_281;
    input [17:0] input_282;
    input [17:0] input_283;
    input [17:0] input_284;
    input [17:0] input_285;
    input [17:0] input_286;
    input [17:0] input_287;
    input [17:0] input_288;
    input [17:0] input_289;
    input [17:0] input_290;
    input [17:0] input_291;
    input [17:0] input_292;
    input [17:0] input_293;
    input [17:0] input_294;
    input [17:0] input_295;
    input [17:0] input_296;
    input [17:0] input_297;
    input [17:0] input_298;
    input [17:0] input_299;
    input [17:0] input_300;
    input [17:0] input_301;
    input [17:0] input_302;
    input [17:0] input_303;
    input [17:0] input_304;
    input [17:0] input_305;
    input [17:0] input_306;
    input [17:0] input_307;
    input [17:0] input_308;
    input [17:0] input_309;
    input [17:0] input_310;
    input [17:0] input_311;
    input [17:0] input_312;
    input [17:0] input_313;
    input [17:0] input_314;
    input [17:0] input_315;
    input [17:0] input_316;
    input [17:0] input_317;
    input [17:0] input_318;
    input [17:0] input_319;
    input [17:0] input_320;
    input [17:0] input_321;
    input [17:0] input_322;
    input [17:0] input_323;
    input [17:0] input_324;
    input [17:0] input_325;
    input [17:0] input_326;
    input [17:0] input_327;
    input [17:0] input_328;
    input [17:0] input_329;
    input [17:0] input_330;
    input [17:0] input_331;
    input [17:0] input_332;
    input [17:0] input_333;
    input [17:0] input_334;
    input [17:0] input_335;
    input [17:0] input_336;
    input [17:0] input_337;
    input [17:0] input_338;
    input [17:0] input_339;
    input [17:0] input_340;
    input [17:0] input_341;
    input [17:0] input_342;
    input [17:0] input_343;
    input [17:0] input_344;
    input [17:0] input_345;
    input [17:0] input_346;
    input [17:0] input_347;
    input [17:0] input_348;
    input [17:0] input_349;
    input [17:0] input_350;
    input [17:0] input_351;
    input [17:0] input_352;
    input [17:0] input_353;
    input [17:0] input_354;
    input [17:0] input_355;
    input [17:0] input_356;
    input [17:0] input_357;
    input [17:0] input_358;
    input [17:0] input_359;
    input [17:0] input_360;
    input [17:0] input_361;
    input [17:0] input_362;
    input [17:0] input_363;
    input [17:0] input_364;
    input [17:0] input_365;
    input [17:0] input_366;
    input [17:0] input_367;
    input [17:0] input_368;
    input [17:0] input_369;
    input [17:0] input_370;
    input [17:0] input_371;
    input [17:0] input_372;
    input [17:0] input_373;
    input [17:0] input_374;
    input [17:0] input_375;
    input [17:0] input_376;
    input [17:0] input_377;
    input [17:0] input_378;
    input [17:0] input_379;
    input [17:0] input_380;
    input [17:0] input_381;
    input [17:0] input_382;
    input [17:0] input_383;
    input [17:0] input_384;
    input [17:0] input_385;
    input [17:0] input_386;
    input [17:0] input_387;
    input [17:0] input_388;
    input [17:0] input_389;
    input [17:0] input_390;
    input [17:0] input_391;
    input [17:0] input_392;
    input [17:0] input_393;
    input [17:0] input_394;
    input [17:0] input_395;
    input [17:0] input_396;
    input [17:0] input_397;
    input [17:0] input_398;
    input [17:0] input_399;
    input [17:0] input_400;
    input [17:0] input_401;
    input [17:0] input_402;
    input [17:0] input_403;
    input [17:0] input_404;
    input [17:0] input_405;
    input [17:0] input_406;
    input [17:0] input_407;
    input [17:0] input_408;
    input [17:0] input_409;
    input [17:0] input_410;
    input [17:0] input_411;
    input [17:0] input_412;
    input [17:0] input_413;
    input [17:0] input_414;
    input [17:0] input_415;
    input [17:0] input_416;
    input [17:0] input_417;
    input [17:0] input_418;
    input [17:0] input_419;
    input [17:0] input_420;
    input [17:0] input_421;
    input [17:0] input_422;
    input [17:0] input_423;
    input [17:0] input_424;
    input [17:0] input_425;
    input [17:0] input_426;
    input [17:0] input_427;
    input [17:0] input_428;
    input [17:0] input_429;
    input [17:0] input_430;
    input [17:0] input_431;
    input [17:0] input_432;
    input [17:0] input_433;
    input [17:0] input_434;
    input [17:0] input_435;
    input [17:0] input_436;
    input [17:0] input_437;
    input [17:0] input_438;
    input [17:0] input_439;
    input [17:0] input_440;
    input [17:0] input_441;
    input [17:0] input_442;
    input [17:0] input_443;
    input [17:0] input_444;
    input [17:0] input_445;
    input [17:0] input_446;
    input [17:0] input_447;
    input [17:0] input_448;
    input [17:0] input_449;
    input [17:0] input_450;
    input [17:0] input_451;
    input [17:0] input_452;
    input [17:0] input_453;
    input [17:0] input_454;
    input [17:0] input_455;
    input [17:0] input_456;
    input [17:0] input_457;
    input [17:0] input_458;
    input [17:0] input_459;
    input [17:0] input_460;
    input [17:0] input_461;
    input [17:0] input_462;
    input [17:0] input_463;
    input [17:0] input_464;
    input [17:0] input_465;
    input [17:0] input_466;
    input [17:0] input_467;
    input [17:0] input_468;
    input [17:0] input_469;
    input [17:0] input_470;
    input [17:0] input_471;
    input [17:0] input_472;
    input [17:0] input_473;
    input [17:0] input_474;
    input [17:0] input_475;
    input [17:0] input_476;
    input [17:0] input_477;
    input [17:0] input_478;
    input [17:0] input_479;
    input [17:0] input_480;
    input [17:0] input_481;
    input [17:0] input_482;
    input [17:0] input_483;
    input [17:0] input_484;
    input [17:0] input_485;
    input [17:0] input_486;
    input [17:0] input_487;
    input [17:0] input_488;
    input [17:0] input_489;
    input [17:0] input_490;
    input [17:0] input_491;
    input [17:0] input_492;
    input [17:0] input_493;
    input [17:0] input_494;
    input [17:0] input_495;
    input [17:0] input_496;
    input [17:0] input_497;
    input [17:0] input_498;
    input [17:0] input_499;
    input [17:0] input_500;
    input [17:0] input_501;
    input [17:0] input_502;
    input [17:0] input_503;
    input [17:0] input_504;
    input [17:0] input_505;
    input [17:0] input_506;
    input [17:0] input_507;
    input [17:0] input_508;
    input [17:0] input_509;
    input [17:0] input_510;
    input [17:0] input_511;
    input [17:0] input_512;
    input [17:0] input_513;
    input [17:0] input_514;
    input [17:0] input_515;
    input [17:0] input_516;
    input [17:0] input_517;
    input [17:0] input_518;
    input [17:0] input_519;
    input [17:0] input_520;
    input [17:0] input_521;
    input [17:0] input_522;
    input [17:0] input_523;
    input [17:0] input_524;
    input [17:0] input_525;
    input [17:0] input_526;
    input [17:0] input_527;
    input [17:0] input_528;
    input [17:0] input_529;
    input [17:0] input_530;
    input [17:0] input_531;
    input [17:0] input_532;
    input [17:0] input_533;
    input [17:0] input_534;
    input [17:0] input_535;
    input [17:0] input_536;
    input [17:0] input_537;
    input [17:0] input_538;
    input [17:0] input_539;
    input [17:0] input_540;
    input [17:0] input_541;
    input [17:0] input_542;
    input [17:0] input_543;
    input [17:0] input_544;
    input [17:0] input_545;
    input [17:0] input_546;
    input [17:0] input_547;
    input [17:0] input_548;
    input [17:0] input_549;
    input [17:0] input_550;
    input [17:0] input_551;
    input [17:0] input_552;
    input [17:0] input_553;
    input [17:0] input_554;
    input [17:0] input_555;
    input [17:0] input_556;
    input [17:0] input_557;
    input [17:0] input_558;
    input [17:0] input_559;
    input [17:0] input_560;
    input [17:0] input_561;
    input [17:0] input_562;
    input [17:0] input_563;
    input [17:0] input_564;
    input [17:0] input_565;
    input [17:0] input_566;
    input [17:0] input_567;
    input [17:0] input_568;
    input [17:0] input_569;
    input [17:0] input_570;
    input [17:0] input_571;
    input [17:0] input_572;
    input [17:0] input_573;
    input [17:0] input_574;
    input [17:0] input_575;
    input [17:0] input_576;
    input [17:0] input_577;
    input [17:0] input_578;
    input [17:0] input_579;
    input [17:0] input_580;
    input [17:0] input_581;
    input [17:0] input_582;
    input [17:0] input_583;
    input [17:0] input_584;
    input [17:0] input_585;
    input [17:0] input_586;
    input [17:0] input_587;
    input [17:0] input_588;
    input [17:0] input_589;
    input [17:0] input_590;
    input [17:0] input_591;
    input [17:0] input_592;
    input [17:0] input_593;
    input [17:0] input_594;
    input [17:0] input_595;
    input [17:0] input_596;
    input [17:0] input_597;
    input [17:0] input_598;
    input [17:0] input_599;
    input [17:0] input_600;
    input [17:0] input_601;
    input [17:0] input_602;
    input [17:0] input_603;
    input [17:0] input_604;
    input [17:0] input_605;
    input [17:0] input_606;
    input [17:0] input_607;
    input [17:0] input_608;
    input [17:0] input_609;
    input [17:0] input_610;
    input [17:0] input_611;
    input [17:0] input_612;
    input [17:0] input_613;
    input [17:0] input_614;
    input [17:0] input_615;
    input [17:0] input_616;
    input [17:0] input_617;
    input [17:0] input_618;
    input [17:0] input_619;
    input [17:0] input_620;
    input [17:0] input_621;
    input [17:0] input_622;
    input [17:0] input_623;
    input [17:0] input_624;
    input [17:0] input_625;
    input [17:0] input_626;
    input [17:0] input_627;
    input [17:0] input_628;
    input [17:0] input_629;
    input [17:0] input_630;
    input [17:0] input_631;
    input [17:0] input_632;
    input [17:0] input_633;
    input [17:0] input_634;
    input [17:0] input_635;
    input [17:0] input_636;
    input [17:0] input_637;
    input [17:0] input_638;
    input [17:0] input_639;
    input [17:0] input_640;
    input [17:0] input_641;
    input [17:0] input_642;
    input [17:0] input_643;
    input [17:0] input_644;
    input [17:0] input_645;
    input [17:0] input_646;
    input [17:0] input_647;
    input [17:0] input_648;
    input [17:0] input_649;
    input [17:0] input_650;
    input [17:0] input_651;
    input [17:0] input_652;
    input [17:0] input_653;
    input [17:0] input_654;
    input [17:0] input_655;
    input [17:0] input_656;
    input [17:0] input_657;
    input [17:0] input_658;
    input [17:0] input_659;
    input [17:0] input_660;
    input [17:0] input_661;
    input [17:0] input_662;
    input [17:0] input_663;
    input [17:0] input_664;
    input [17:0] input_665;
    input [17:0] input_666;
    input [17:0] input_667;
    input [17:0] input_668;
    input [17:0] input_669;
    input [17:0] input_670;
    input [17:0] input_671;
    input [17:0] input_672;
    input [17:0] input_673;
    input [17:0] input_674;
    input [17:0] input_675;
    input [17:0] input_676;
    input [17:0] input_677;
    input [17:0] input_678;
    input [17:0] input_679;
    input [17:0] input_680;
    input [17:0] input_681;
    input [17:0] input_682;
    input [17:0] input_683;
    input [17:0] input_684;
    input [17:0] input_685;
    input [17:0] input_686;
    input [17:0] input_687;
    input [17:0] input_688;
    input [17:0] input_689;
    input [17:0] input_690;
    input [17:0] input_691;
    input [17:0] input_692;
    input [17:0] input_693;
    input [17:0] input_694;
    input [17:0] input_695;
    input [17:0] input_696;
    input [17:0] input_697;
    input [17:0] input_698;
    input [17:0] input_699;
    input [17:0] input_700;
    input [17:0] input_701;
    input [17:0] input_702;
    input [17:0] input_703;
    input [17:0] input_704;
    input [17:0] input_705;
    input [17:0] input_706;
    input [17:0] input_707;
    input [17:0] input_708;
    input [17:0] input_709;
    input [17:0] input_710;
    input [17:0] input_711;
    input [17:0] input_712;
    input [17:0] input_713;
    input [17:0] input_714;
    input [17:0] input_715;
    input [17:0] input_716;
    input [17:0] input_717;
    input [17:0] input_718;
    input [17:0] input_719;
    input [17:0] input_720;
    input [17:0] input_721;
    input [17:0] input_722;
    input [17:0] input_723;
    input [17:0] input_724;
    input [17:0] input_725;
    input [17:0] input_726;
    input [17:0] input_727;
    input [17:0] input_728;
    input [17:0] input_729;
    input [17:0] input_730;
    input [17:0] input_731;
    input [17:0] input_732;
    input [17:0] input_733;
    input [17:0] input_734;
    input [17:0] input_735;
    input [17:0] input_736;
    input [17:0] input_737;
    input [17:0] input_738;
    input [17:0] input_739;
    input [17:0] input_740;
    input [17:0] input_741;
    input [17:0] input_742;
    input [17:0] input_743;
    input [17:0] input_744;
    input [17:0] input_745;
    input [17:0] input_746;
    input [17:0] input_747;
    input [17:0] input_748;
    input [17:0] input_749;
    input [17:0] input_750;
    input [17:0] input_751;
    input [17:0] input_752;
    input [17:0] input_753;
    input [17:0] input_754;
    input [17:0] input_755;
    input [17:0] input_756;
    input [17:0] input_757;
    input [17:0] input_758;
    input [17:0] input_759;
    input [17:0] input_760;
    input [17:0] input_761;
    input [17:0] input_762;
    input [17:0] input_763;
    input [17:0] input_764;
    input [17:0] input_765;
    input [17:0] input_766;
    input [17:0] input_767;
    input [17:0] input_768;
    input [17:0] input_769;
    input [17:0] input_770;
    input [17:0] input_771;
    input [17:0] input_772;
    input [17:0] input_773;
    input [17:0] input_774;
    input [17:0] input_775;
    input [17:0] input_776;
    input [17:0] input_777;
    input [17:0] input_778;
    input [17:0] input_779;
    input [17:0] input_780;
    input [17:0] input_781;
    input [17:0] input_782;
    input [17:0] input_783;
    input [9:0] sel;
    reg [17:0] result;
  begin
    case (sel)
      10'b0000000000 : begin
        result = input_0;
      end
      10'b0000000001 : begin
        result = input_1;
      end
      10'b0000000010 : begin
        result = input_2;
      end
      10'b0000000011 : begin
        result = input_3;
      end
      10'b0000000100 : begin
        result = input_4;
      end
      10'b0000000101 : begin
        result = input_5;
      end
      10'b0000000110 : begin
        result = input_6;
      end
      10'b0000000111 : begin
        result = input_7;
      end
      10'b0000001000 : begin
        result = input_8;
      end
      10'b0000001001 : begin
        result = input_9;
      end
      10'b0000001010 : begin
        result = input_10;
      end
      10'b0000001011 : begin
        result = input_11;
      end
      10'b0000001100 : begin
        result = input_12;
      end
      10'b0000001101 : begin
        result = input_13;
      end
      10'b0000001110 : begin
        result = input_14;
      end
      10'b0000001111 : begin
        result = input_15;
      end
      10'b0000010000 : begin
        result = input_16;
      end
      10'b0000010001 : begin
        result = input_17;
      end
      10'b0000010010 : begin
        result = input_18;
      end
      10'b0000010011 : begin
        result = input_19;
      end
      10'b0000010100 : begin
        result = input_20;
      end
      10'b0000010101 : begin
        result = input_21;
      end
      10'b0000010110 : begin
        result = input_22;
      end
      10'b0000010111 : begin
        result = input_23;
      end
      10'b0000011000 : begin
        result = input_24;
      end
      10'b0000011001 : begin
        result = input_25;
      end
      10'b0000011010 : begin
        result = input_26;
      end
      10'b0000011011 : begin
        result = input_27;
      end
      10'b0000011100 : begin
        result = input_28;
      end
      10'b0000011101 : begin
        result = input_29;
      end
      10'b0000011110 : begin
        result = input_30;
      end
      10'b0000011111 : begin
        result = input_31;
      end
      10'b0000100000 : begin
        result = input_32;
      end
      10'b0000100001 : begin
        result = input_33;
      end
      10'b0000100010 : begin
        result = input_34;
      end
      10'b0000100011 : begin
        result = input_35;
      end
      10'b0000100100 : begin
        result = input_36;
      end
      10'b0000100101 : begin
        result = input_37;
      end
      10'b0000100110 : begin
        result = input_38;
      end
      10'b0000100111 : begin
        result = input_39;
      end
      10'b0000101000 : begin
        result = input_40;
      end
      10'b0000101001 : begin
        result = input_41;
      end
      10'b0000101010 : begin
        result = input_42;
      end
      10'b0000101011 : begin
        result = input_43;
      end
      10'b0000101100 : begin
        result = input_44;
      end
      10'b0000101101 : begin
        result = input_45;
      end
      10'b0000101110 : begin
        result = input_46;
      end
      10'b0000101111 : begin
        result = input_47;
      end
      10'b0000110000 : begin
        result = input_48;
      end
      10'b0000110001 : begin
        result = input_49;
      end
      10'b0000110010 : begin
        result = input_50;
      end
      10'b0000110011 : begin
        result = input_51;
      end
      10'b0000110100 : begin
        result = input_52;
      end
      10'b0000110101 : begin
        result = input_53;
      end
      10'b0000110110 : begin
        result = input_54;
      end
      10'b0000110111 : begin
        result = input_55;
      end
      10'b0000111000 : begin
        result = input_56;
      end
      10'b0000111001 : begin
        result = input_57;
      end
      10'b0000111010 : begin
        result = input_58;
      end
      10'b0000111011 : begin
        result = input_59;
      end
      10'b0000111100 : begin
        result = input_60;
      end
      10'b0000111101 : begin
        result = input_61;
      end
      10'b0000111110 : begin
        result = input_62;
      end
      10'b0000111111 : begin
        result = input_63;
      end
      10'b0001000000 : begin
        result = input_64;
      end
      10'b0001000001 : begin
        result = input_65;
      end
      10'b0001000010 : begin
        result = input_66;
      end
      10'b0001000011 : begin
        result = input_67;
      end
      10'b0001000100 : begin
        result = input_68;
      end
      10'b0001000101 : begin
        result = input_69;
      end
      10'b0001000110 : begin
        result = input_70;
      end
      10'b0001000111 : begin
        result = input_71;
      end
      10'b0001001000 : begin
        result = input_72;
      end
      10'b0001001001 : begin
        result = input_73;
      end
      10'b0001001010 : begin
        result = input_74;
      end
      10'b0001001011 : begin
        result = input_75;
      end
      10'b0001001100 : begin
        result = input_76;
      end
      10'b0001001101 : begin
        result = input_77;
      end
      10'b0001001110 : begin
        result = input_78;
      end
      10'b0001001111 : begin
        result = input_79;
      end
      10'b0001010000 : begin
        result = input_80;
      end
      10'b0001010001 : begin
        result = input_81;
      end
      10'b0001010010 : begin
        result = input_82;
      end
      10'b0001010011 : begin
        result = input_83;
      end
      10'b0001010100 : begin
        result = input_84;
      end
      10'b0001010101 : begin
        result = input_85;
      end
      10'b0001010110 : begin
        result = input_86;
      end
      10'b0001010111 : begin
        result = input_87;
      end
      10'b0001011000 : begin
        result = input_88;
      end
      10'b0001011001 : begin
        result = input_89;
      end
      10'b0001011010 : begin
        result = input_90;
      end
      10'b0001011011 : begin
        result = input_91;
      end
      10'b0001011100 : begin
        result = input_92;
      end
      10'b0001011101 : begin
        result = input_93;
      end
      10'b0001011110 : begin
        result = input_94;
      end
      10'b0001011111 : begin
        result = input_95;
      end
      10'b0001100000 : begin
        result = input_96;
      end
      10'b0001100001 : begin
        result = input_97;
      end
      10'b0001100010 : begin
        result = input_98;
      end
      10'b0001100011 : begin
        result = input_99;
      end
      10'b0001100100 : begin
        result = input_100;
      end
      10'b0001100101 : begin
        result = input_101;
      end
      10'b0001100110 : begin
        result = input_102;
      end
      10'b0001100111 : begin
        result = input_103;
      end
      10'b0001101000 : begin
        result = input_104;
      end
      10'b0001101001 : begin
        result = input_105;
      end
      10'b0001101010 : begin
        result = input_106;
      end
      10'b0001101011 : begin
        result = input_107;
      end
      10'b0001101100 : begin
        result = input_108;
      end
      10'b0001101101 : begin
        result = input_109;
      end
      10'b0001101110 : begin
        result = input_110;
      end
      10'b0001101111 : begin
        result = input_111;
      end
      10'b0001110000 : begin
        result = input_112;
      end
      10'b0001110001 : begin
        result = input_113;
      end
      10'b0001110010 : begin
        result = input_114;
      end
      10'b0001110011 : begin
        result = input_115;
      end
      10'b0001110100 : begin
        result = input_116;
      end
      10'b0001110101 : begin
        result = input_117;
      end
      10'b0001110110 : begin
        result = input_118;
      end
      10'b0001110111 : begin
        result = input_119;
      end
      10'b0001111000 : begin
        result = input_120;
      end
      10'b0001111001 : begin
        result = input_121;
      end
      10'b0001111010 : begin
        result = input_122;
      end
      10'b0001111011 : begin
        result = input_123;
      end
      10'b0001111100 : begin
        result = input_124;
      end
      10'b0001111101 : begin
        result = input_125;
      end
      10'b0001111110 : begin
        result = input_126;
      end
      10'b0001111111 : begin
        result = input_127;
      end
      10'b0010000000 : begin
        result = input_128;
      end
      10'b0010000001 : begin
        result = input_129;
      end
      10'b0010000010 : begin
        result = input_130;
      end
      10'b0010000011 : begin
        result = input_131;
      end
      10'b0010000100 : begin
        result = input_132;
      end
      10'b0010000101 : begin
        result = input_133;
      end
      10'b0010000110 : begin
        result = input_134;
      end
      10'b0010000111 : begin
        result = input_135;
      end
      10'b0010001000 : begin
        result = input_136;
      end
      10'b0010001001 : begin
        result = input_137;
      end
      10'b0010001010 : begin
        result = input_138;
      end
      10'b0010001011 : begin
        result = input_139;
      end
      10'b0010001100 : begin
        result = input_140;
      end
      10'b0010001101 : begin
        result = input_141;
      end
      10'b0010001110 : begin
        result = input_142;
      end
      10'b0010001111 : begin
        result = input_143;
      end
      10'b0010010000 : begin
        result = input_144;
      end
      10'b0010010001 : begin
        result = input_145;
      end
      10'b0010010010 : begin
        result = input_146;
      end
      10'b0010010011 : begin
        result = input_147;
      end
      10'b0010010100 : begin
        result = input_148;
      end
      10'b0010010101 : begin
        result = input_149;
      end
      10'b0010010110 : begin
        result = input_150;
      end
      10'b0010010111 : begin
        result = input_151;
      end
      10'b0010011000 : begin
        result = input_152;
      end
      10'b0010011001 : begin
        result = input_153;
      end
      10'b0010011010 : begin
        result = input_154;
      end
      10'b0010011011 : begin
        result = input_155;
      end
      10'b0010011100 : begin
        result = input_156;
      end
      10'b0010011101 : begin
        result = input_157;
      end
      10'b0010011110 : begin
        result = input_158;
      end
      10'b0010011111 : begin
        result = input_159;
      end
      10'b0010100000 : begin
        result = input_160;
      end
      10'b0010100001 : begin
        result = input_161;
      end
      10'b0010100010 : begin
        result = input_162;
      end
      10'b0010100011 : begin
        result = input_163;
      end
      10'b0010100100 : begin
        result = input_164;
      end
      10'b0010100101 : begin
        result = input_165;
      end
      10'b0010100110 : begin
        result = input_166;
      end
      10'b0010100111 : begin
        result = input_167;
      end
      10'b0010101000 : begin
        result = input_168;
      end
      10'b0010101001 : begin
        result = input_169;
      end
      10'b0010101010 : begin
        result = input_170;
      end
      10'b0010101011 : begin
        result = input_171;
      end
      10'b0010101100 : begin
        result = input_172;
      end
      10'b0010101101 : begin
        result = input_173;
      end
      10'b0010101110 : begin
        result = input_174;
      end
      10'b0010101111 : begin
        result = input_175;
      end
      10'b0010110000 : begin
        result = input_176;
      end
      10'b0010110001 : begin
        result = input_177;
      end
      10'b0010110010 : begin
        result = input_178;
      end
      10'b0010110011 : begin
        result = input_179;
      end
      10'b0010110100 : begin
        result = input_180;
      end
      10'b0010110101 : begin
        result = input_181;
      end
      10'b0010110110 : begin
        result = input_182;
      end
      10'b0010110111 : begin
        result = input_183;
      end
      10'b0010111000 : begin
        result = input_184;
      end
      10'b0010111001 : begin
        result = input_185;
      end
      10'b0010111010 : begin
        result = input_186;
      end
      10'b0010111011 : begin
        result = input_187;
      end
      10'b0010111100 : begin
        result = input_188;
      end
      10'b0010111101 : begin
        result = input_189;
      end
      10'b0010111110 : begin
        result = input_190;
      end
      10'b0010111111 : begin
        result = input_191;
      end
      10'b0011000000 : begin
        result = input_192;
      end
      10'b0011000001 : begin
        result = input_193;
      end
      10'b0011000010 : begin
        result = input_194;
      end
      10'b0011000011 : begin
        result = input_195;
      end
      10'b0011000100 : begin
        result = input_196;
      end
      10'b0011000101 : begin
        result = input_197;
      end
      10'b0011000110 : begin
        result = input_198;
      end
      10'b0011000111 : begin
        result = input_199;
      end
      10'b0011001000 : begin
        result = input_200;
      end
      10'b0011001001 : begin
        result = input_201;
      end
      10'b0011001010 : begin
        result = input_202;
      end
      10'b0011001011 : begin
        result = input_203;
      end
      10'b0011001100 : begin
        result = input_204;
      end
      10'b0011001101 : begin
        result = input_205;
      end
      10'b0011001110 : begin
        result = input_206;
      end
      10'b0011001111 : begin
        result = input_207;
      end
      10'b0011010000 : begin
        result = input_208;
      end
      10'b0011010001 : begin
        result = input_209;
      end
      10'b0011010010 : begin
        result = input_210;
      end
      10'b0011010011 : begin
        result = input_211;
      end
      10'b0011010100 : begin
        result = input_212;
      end
      10'b0011010101 : begin
        result = input_213;
      end
      10'b0011010110 : begin
        result = input_214;
      end
      10'b0011010111 : begin
        result = input_215;
      end
      10'b0011011000 : begin
        result = input_216;
      end
      10'b0011011001 : begin
        result = input_217;
      end
      10'b0011011010 : begin
        result = input_218;
      end
      10'b0011011011 : begin
        result = input_219;
      end
      10'b0011011100 : begin
        result = input_220;
      end
      10'b0011011101 : begin
        result = input_221;
      end
      10'b0011011110 : begin
        result = input_222;
      end
      10'b0011011111 : begin
        result = input_223;
      end
      10'b0011100000 : begin
        result = input_224;
      end
      10'b0011100001 : begin
        result = input_225;
      end
      10'b0011100010 : begin
        result = input_226;
      end
      10'b0011100011 : begin
        result = input_227;
      end
      10'b0011100100 : begin
        result = input_228;
      end
      10'b0011100101 : begin
        result = input_229;
      end
      10'b0011100110 : begin
        result = input_230;
      end
      10'b0011100111 : begin
        result = input_231;
      end
      10'b0011101000 : begin
        result = input_232;
      end
      10'b0011101001 : begin
        result = input_233;
      end
      10'b0011101010 : begin
        result = input_234;
      end
      10'b0011101011 : begin
        result = input_235;
      end
      10'b0011101100 : begin
        result = input_236;
      end
      10'b0011101101 : begin
        result = input_237;
      end
      10'b0011101110 : begin
        result = input_238;
      end
      10'b0011101111 : begin
        result = input_239;
      end
      10'b0011110000 : begin
        result = input_240;
      end
      10'b0011110001 : begin
        result = input_241;
      end
      10'b0011110010 : begin
        result = input_242;
      end
      10'b0011110011 : begin
        result = input_243;
      end
      10'b0011110100 : begin
        result = input_244;
      end
      10'b0011110101 : begin
        result = input_245;
      end
      10'b0011110110 : begin
        result = input_246;
      end
      10'b0011110111 : begin
        result = input_247;
      end
      10'b0011111000 : begin
        result = input_248;
      end
      10'b0011111001 : begin
        result = input_249;
      end
      10'b0011111010 : begin
        result = input_250;
      end
      10'b0011111011 : begin
        result = input_251;
      end
      10'b0011111100 : begin
        result = input_252;
      end
      10'b0011111101 : begin
        result = input_253;
      end
      10'b0011111110 : begin
        result = input_254;
      end
      10'b0011111111 : begin
        result = input_255;
      end
      10'b0100000000 : begin
        result = input_256;
      end
      10'b0100000001 : begin
        result = input_257;
      end
      10'b0100000010 : begin
        result = input_258;
      end
      10'b0100000011 : begin
        result = input_259;
      end
      10'b0100000100 : begin
        result = input_260;
      end
      10'b0100000101 : begin
        result = input_261;
      end
      10'b0100000110 : begin
        result = input_262;
      end
      10'b0100000111 : begin
        result = input_263;
      end
      10'b0100001000 : begin
        result = input_264;
      end
      10'b0100001001 : begin
        result = input_265;
      end
      10'b0100001010 : begin
        result = input_266;
      end
      10'b0100001011 : begin
        result = input_267;
      end
      10'b0100001100 : begin
        result = input_268;
      end
      10'b0100001101 : begin
        result = input_269;
      end
      10'b0100001110 : begin
        result = input_270;
      end
      10'b0100001111 : begin
        result = input_271;
      end
      10'b0100010000 : begin
        result = input_272;
      end
      10'b0100010001 : begin
        result = input_273;
      end
      10'b0100010010 : begin
        result = input_274;
      end
      10'b0100010011 : begin
        result = input_275;
      end
      10'b0100010100 : begin
        result = input_276;
      end
      10'b0100010101 : begin
        result = input_277;
      end
      10'b0100010110 : begin
        result = input_278;
      end
      10'b0100010111 : begin
        result = input_279;
      end
      10'b0100011000 : begin
        result = input_280;
      end
      10'b0100011001 : begin
        result = input_281;
      end
      10'b0100011010 : begin
        result = input_282;
      end
      10'b0100011011 : begin
        result = input_283;
      end
      10'b0100011100 : begin
        result = input_284;
      end
      10'b0100011101 : begin
        result = input_285;
      end
      10'b0100011110 : begin
        result = input_286;
      end
      10'b0100011111 : begin
        result = input_287;
      end
      10'b0100100000 : begin
        result = input_288;
      end
      10'b0100100001 : begin
        result = input_289;
      end
      10'b0100100010 : begin
        result = input_290;
      end
      10'b0100100011 : begin
        result = input_291;
      end
      10'b0100100100 : begin
        result = input_292;
      end
      10'b0100100101 : begin
        result = input_293;
      end
      10'b0100100110 : begin
        result = input_294;
      end
      10'b0100100111 : begin
        result = input_295;
      end
      10'b0100101000 : begin
        result = input_296;
      end
      10'b0100101001 : begin
        result = input_297;
      end
      10'b0100101010 : begin
        result = input_298;
      end
      10'b0100101011 : begin
        result = input_299;
      end
      10'b0100101100 : begin
        result = input_300;
      end
      10'b0100101101 : begin
        result = input_301;
      end
      10'b0100101110 : begin
        result = input_302;
      end
      10'b0100101111 : begin
        result = input_303;
      end
      10'b0100110000 : begin
        result = input_304;
      end
      10'b0100110001 : begin
        result = input_305;
      end
      10'b0100110010 : begin
        result = input_306;
      end
      10'b0100110011 : begin
        result = input_307;
      end
      10'b0100110100 : begin
        result = input_308;
      end
      10'b0100110101 : begin
        result = input_309;
      end
      10'b0100110110 : begin
        result = input_310;
      end
      10'b0100110111 : begin
        result = input_311;
      end
      10'b0100111000 : begin
        result = input_312;
      end
      10'b0100111001 : begin
        result = input_313;
      end
      10'b0100111010 : begin
        result = input_314;
      end
      10'b0100111011 : begin
        result = input_315;
      end
      10'b0100111100 : begin
        result = input_316;
      end
      10'b0100111101 : begin
        result = input_317;
      end
      10'b0100111110 : begin
        result = input_318;
      end
      10'b0100111111 : begin
        result = input_319;
      end
      10'b0101000000 : begin
        result = input_320;
      end
      10'b0101000001 : begin
        result = input_321;
      end
      10'b0101000010 : begin
        result = input_322;
      end
      10'b0101000011 : begin
        result = input_323;
      end
      10'b0101000100 : begin
        result = input_324;
      end
      10'b0101000101 : begin
        result = input_325;
      end
      10'b0101000110 : begin
        result = input_326;
      end
      10'b0101000111 : begin
        result = input_327;
      end
      10'b0101001000 : begin
        result = input_328;
      end
      10'b0101001001 : begin
        result = input_329;
      end
      10'b0101001010 : begin
        result = input_330;
      end
      10'b0101001011 : begin
        result = input_331;
      end
      10'b0101001100 : begin
        result = input_332;
      end
      10'b0101001101 : begin
        result = input_333;
      end
      10'b0101001110 : begin
        result = input_334;
      end
      10'b0101001111 : begin
        result = input_335;
      end
      10'b0101010000 : begin
        result = input_336;
      end
      10'b0101010001 : begin
        result = input_337;
      end
      10'b0101010010 : begin
        result = input_338;
      end
      10'b0101010011 : begin
        result = input_339;
      end
      10'b0101010100 : begin
        result = input_340;
      end
      10'b0101010101 : begin
        result = input_341;
      end
      10'b0101010110 : begin
        result = input_342;
      end
      10'b0101010111 : begin
        result = input_343;
      end
      10'b0101011000 : begin
        result = input_344;
      end
      10'b0101011001 : begin
        result = input_345;
      end
      10'b0101011010 : begin
        result = input_346;
      end
      10'b0101011011 : begin
        result = input_347;
      end
      10'b0101011100 : begin
        result = input_348;
      end
      10'b0101011101 : begin
        result = input_349;
      end
      10'b0101011110 : begin
        result = input_350;
      end
      10'b0101011111 : begin
        result = input_351;
      end
      10'b0101100000 : begin
        result = input_352;
      end
      10'b0101100001 : begin
        result = input_353;
      end
      10'b0101100010 : begin
        result = input_354;
      end
      10'b0101100011 : begin
        result = input_355;
      end
      10'b0101100100 : begin
        result = input_356;
      end
      10'b0101100101 : begin
        result = input_357;
      end
      10'b0101100110 : begin
        result = input_358;
      end
      10'b0101100111 : begin
        result = input_359;
      end
      10'b0101101000 : begin
        result = input_360;
      end
      10'b0101101001 : begin
        result = input_361;
      end
      10'b0101101010 : begin
        result = input_362;
      end
      10'b0101101011 : begin
        result = input_363;
      end
      10'b0101101100 : begin
        result = input_364;
      end
      10'b0101101101 : begin
        result = input_365;
      end
      10'b0101101110 : begin
        result = input_366;
      end
      10'b0101101111 : begin
        result = input_367;
      end
      10'b0101110000 : begin
        result = input_368;
      end
      10'b0101110001 : begin
        result = input_369;
      end
      10'b0101110010 : begin
        result = input_370;
      end
      10'b0101110011 : begin
        result = input_371;
      end
      10'b0101110100 : begin
        result = input_372;
      end
      10'b0101110101 : begin
        result = input_373;
      end
      10'b0101110110 : begin
        result = input_374;
      end
      10'b0101110111 : begin
        result = input_375;
      end
      10'b0101111000 : begin
        result = input_376;
      end
      10'b0101111001 : begin
        result = input_377;
      end
      10'b0101111010 : begin
        result = input_378;
      end
      10'b0101111011 : begin
        result = input_379;
      end
      10'b0101111100 : begin
        result = input_380;
      end
      10'b0101111101 : begin
        result = input_381;
      end
      10'b0101111110 : begin
        result = input_382;
      end
      10'b0101111111 : begin
        result = input_383;
      end
      10'b0110000000 : begin
        result = input_384;
      end
      10'b0110000001 : begin
        result = input_385;
      end
      10'b0110000010 : begin
        result = input_386;
      end
      10'b0110000011 : begin
        result = input_387;
      end
      10'b0110000100 : begin
        result = input_388;
      end
      10'b0110000101 : begin
        result = input_389;
      end
      10'b0110000110 : begin
        result = input_390;
      end
      10'b0110000111 : begin
        result = input_391;
      end
      10'b0110001000 : begin
        result = input_392;
      end
      10'b0110001001 : begin
        result = input_393;
      end
      10'b0110001010 : begin
        result = input_394;
      end
      10'b0110001011 : begin
        result = input_395;
      end
      10'b0110001100 : begin
        result = input_396;
      end
      10'b0110001101 : begin
        result = input_397;
      end
      10'b0110001110 : begin
        result = input_398;
      end
      10'b0110001111 : begin
        result = input_399;
      end
      10'b0110010000 : begin
        result = input_400;
      end
      10'b0110010001 : begin
        result = input_401;
      end
      10'b0110010010 : begin
        result = input_402;
      end
      10'b0110010011 : begin
        result = input_403;
      end
      10'b0110010100 : begin
        result = input_404;
      end
      10'b0110010101 : begin
        result = input_405;
      end
      10'b0110010110 : begin
        result = input_406;
      end
      10'b0110010111 : begin
        result = input_407;
      end
      10'b0110011000 : begin
        result = input_408;
      end
      10'b0110011001 : begin
        result = input_409;
      end
      10'b0110011010 : begin
        result = input_410;
      end
      10'b0110011011 : begin
        result = input_411;
      end
      10'b0110011100 : begin
        result = input_412;
      end
      10'b0110011101 : begin
        result = input_413;
      end
      10'b0110011110 : begin
        result = input_414;
      end
      10'b0110011111 : begin
        result = input_415;
      end
      10'b0110100000 : begin
        result = input_416;
      end
      10'b0110100001 : begin
        result = input_417;
      end
      10'b0110100010 : begin
        result = input_418;
      end
      10'b0110100011 : begin
        result = input_419;
      end
      10'b0110100100 : begin
        result = input_420;
      end
      10'b0110100101 : begin
        result = input_421;
      end
      10'b0110100110 : begin
        result = input_422;
      end
      10'b0110100111 : begin
        result = input_423;
      end
      10'b0110101000 : begin
        result = input_424;
      end
      10'b0110101001 : begin
        result = input_425;
      end
      10'b0110101010 : begin
        result = input_426;
      end
      10'b0110101011 : begin
        result = input_427;
      end
      10'b0110101100 : begin
        result = input_428;
      end
      10'b0110101101 : begin
        result = input_429;
      end
      10'b0110101110 : begin
        result = input_430;
      end
      10'b0110101111 : begin
        result = input_431;
      end
      10'b0110110000 : begin
        result = input_432;
      end
      10'b0110110001 : begin
        result = input_433;
      end
      10'b0110110010 : begin
        result = input_434;
      end
      10'b0110110011 : begin
        result = input_435;
      end
      10'b0110110100 : begin
        result = input_436;
      end
      10'b0110110101 : begin
        result = input_437;
      end
      10'b0110110110 : begin
        result = input_438;
      end
      10'b0110110111 : begin
        result = input_439;
      end
      10'b0110111000 : begin
        result = input_440;
      end
      10'b0110111001 : begin
        result = input_441;
      end
      10'b0110111010 : begin
        result = input_442;
      end
      10'b0110111011 : begin
        result = input_443;
      end
      10'b0110111100 : begin
        result = input_444;
      end
      10'b0110111101 : begin
        result = input_445;
      end
      10'b0110111110 : begin
        result = input_446;
      end
      10'b0110111111 : begin
        result = input_447;
      end
      10'b0111000000 : begin
        result = input_448;
      end
      10'b0111000001 : begin
        result = input_449;
      end
      10'b0111000010 : begin
        result = input_450;
      end
      10'b0111000011 : begin
        result = input_451;
      end
      10'b0111000100 : begin
        result = input_452;
      end
      10'b0111000101 : begin
        result = input_453;
      end
      10'b0111000110 : begin
        result = input_454;
      end
      10'b0111000111 : begin
        result = input_455;
      end
      10'b0111001000 : begin
        result = input_456;
      end
      10'b0111001001 : begin
        result = input_457;
      end
      10'b0111001010 : begin
        result = input_458;
      end
      10'b0111001011 : begin
        result = input_459;
      end
      10'b0111001100 : begin
        result = input_460;
      end
      10'b0111001101 : begin
        result = input_461;
      end
      10'b0111001110 : begin
        result = input_462;
      end
      10'b0111001111 : begin
        result = input_463;
      end
      10'b0111010000 : begin
        result = input_464;
      end
      10'b0111010001 : begin
        result = input_465;
      end
      10'b0111010010 : begin
        result = input_466;
      end
      10'b0111010011 : begin
        result = input_467;
      end
      10'b0111010100 : begin
        result = input_468;
      end
      10'b0111010101 : begin
        result = input_469;
      end
      10'b0111010110 : begin
        result = input_470;
      end
      10'b0111010111 : begin
        result = input_471;
      end
      10'b0111011000 : begin
        result = input_472;
      end
      10'b0111011001 : begin
        result = input_473;
      end
      10'b0111011010 : begin
        result = input_474;
      end
      10'b0111011011 : begin
        result = input_475;
      end
      10'b0111011100 : begin
        result = input_476;
      end
      10'b0111011101 : begin
        result = input_477;
      end
      10'b0111011110 : begin
        result = input_478;
      end
      10'b0111011111 : begin
        result = input_479;
      end
      10'b0111100000 : begin
        result = input_480;
      end
      10'b0111100001 : begin
        result = input_481;
      end
      10'b0111100010 : begin
        result = input_482;
      end
      10'b0111100011 : begin
        result = input_483;
      end
      10'b0111100100 : begin
        result = input_484;
      end
      10'b0111100101 : begin
        result = input_485;
      end
      10'b0111100110 : begin
        result = input_486;
      end
      10'b0111100111 : begin
        result = input_487;
      end
      10'b0111101000 : begin
        result = input_488;
      end
      10'b0111101001 : begin
        result = input_489;
      end
      10'b0111101010 : begin
        result = input_490;
      end
      10'b0111101011 : begin
        result = input_491;
      end
      10'b0111101100 : begin
        result = input_492;
      end
      10'b0111101101 : begin
        result = input_493;
      end
      10'b0111101110 : begin
        result = input_494;
      end
      10'b0111101111 : begin
        result = input_495;
      end
      10'b0111110000 : begin
        result = input_496;
      end
      10'b0111110001 : begin
        result = input_497;
      end
      10'b0111110010 : begin
        result = input_498;
      end
      10'b0111110011 : begin
        result = input_499;
      end
      10'b0111110100 : begin
        result = input_500;
      end
      10'b0111110101 : begin
        result = input_501;
      end
      10'b0111110110 : begin
        result = input_502;
      end
      10'b0111110111 : begin
        result = input_503;
      end
      10'b0111111000 : begin
        result = input_504;
      end
      10'b0111111001 : begin
        result = input_505;
      end
      10'b0111111010 : begin
        result = input_506;
      end
      10'b0111111011 : begin
        result = input_507;
      end
      10'b0111111100 : begin
        result = input_508;
      end
      10'b0111111101 : begin
        result = input_509;
      end
      10'b0111111110 : begin
        result = input_510;
      end
      10'b0111111111 : begin
        result = input_511;
      end
      10'b1000000000 : begin
        result = input_512;
      end
      10'b1000000001 : begin
        result = input_513;
      end
      10'b1000000010 : begin
        result = input_514;
      end
      10'b1000000011 : begin
        result = input_515;
      end
      10'b1000000100 : begin
        result = input_516;
      end
      10'b1000000101 : begin
        result = input_517;
      end
      10'b1000000110 : begin
        result = input_518;
      end
      10'b1000000111 : begin
        result = input_519;
      end
      10'b1000001000 : begin
        result = input_520;
      end
      10'b1000001001 : begin
        result = input_521;
      end
      10'b1000001010 : begin
        result = input_522;
      end
      10'b1000001011 : begin
        result = input_523;
      end
      10'b1000001100 : begin
        result = input_524;
      end
      10'b1000001101 : begin
        result = input_525;
      end
      10'b1000001110 : begin
        result = input_526;
      end
      10'b1000001111 : begin
        result = input_527;
      end
      10'b1000010000 : begin
        result = input_528;
      end
      10'b1000010001 : begin
        result = input_529;
      end
      10'b1000010010 : begin
        result = input_530;
      end
      10'b1000010011 : begin
        result = input_531;
      end
      10'b1000010100 : begin
        result = input_532;
      end
      10'b1000010101 : begin
        result = input_533;
      end
      10'b1000010110 : begin
        result = input_534;
      end
      10'b1000010111 : begin
        result = input_535;
      end
      10'b1000011000 : begin
        result = input_536;
      end
      10'b1000011001 : begin
        result = input_537;
      end
      10'b1000011010 : begin
        result = input_538;
      end
      10'b1000011011 : begin
        result = input_539;
      end
      10'b1000011100 : begin
        result = input_540;
      end
      10'b1000011101 : begin
        result = input_541;
      end
      10'b1000011110 : begin
        result = input_542;
      end
      10'b1000011111 : begin
        result = input_543;
      end
      10'b1000100000 : begin
        result = input_544;
      end
      10'b1000100001 : begin
        result = input_545;
      end
      10'b1000100010 : begin
        result = input_546;
      end
      10'b1000100011 : begin
        result = input_547;
      end
      10'b1000100100 : begin
        result = input_548;
      end
      10'b1000100101 : begin
        result = input_549;
      end
      10'b1000100110 : begin
        result = input_550;
      end
      10'b1000100111 : begin
        result = input_551;
      end
      10'b1000101000 : begin
        result = input_552;
      end
      10'b1000101001 : begin
        result = input_553;
      end
      10'b1000101010 : begin
        result = input_554;
      end
      10'b1000101011 : begin
        result = input_555;
      end
      10'b1000101100 : begin
        result = input_556;
      end
      10'b1000101101 : begin
        result = input_557;
      end
      10'b1000101110 : begin
        result = input_558;
      end
      10'b1000101111 : begin
        result = input_559;
      end
      10'b1000110000 : begin
        result = input_560;
      end
      10'b1000110001 : begin
        result = input_561;
      end
      10'b1000110010 : begin
        result = input_562;
      end
      10'b1000110011 : begin
        result = input_563;
      end
      10'b1000110100 : begin
        result = input_564;
      end
      10'b1000110101 : begin
        result = input_565;
      end
      10'b1000110110 : begin
        result = input_566;
      end
      10'b1000110111 : begin
        result = input_567;
      end
      10'b1000111000 : begin
        result = input_568;
      end
      10'b1000111001 : begin
        result = input_569;
      end
      10'b1000111010 : begin
        result = input_570;
      end
      10'b1000111011 : begin
        result = input_571;
      end
      10'b1000111100 : begin
        result = input_572;
      end
      10'b1000111101 : begin
        result = input_573;
      end
      10'b1000111110 : begin
        result = input_574;
      end
      10'b1000111111 : begin
        result = input_575;
      end
      10'b1001000000 : begin
        result = input_576;
      end
      10'b1001000001 : begin
        result = input_577;
      end
      10'b1001000010 : begin
        result = input_578;
      end
      10'b1001000011 : begin
        result = input_579;
      end
      10'b1001000100 : begin
        result = input_580;
      end
      10'b1001000101 : begin
        result = input_581;
      end
      10'b1001000110 : begin
        result = input_582;
      end
      10'b1001000111 : begin
        result = input_583;
      end
      10'b1001001000 : begin
        result = input_584;
      end
      10'b1001001001 : begin
        result = input_585;
      end
      10'b1001001010 : begin
        result = input_586;
      end
      10'b1001001011 : begin
        result = input_587;
      end
      10'b1001001100 : begin
        result = input_588;
      end
      10'b1001001101 : begin
        result = input_589;
      end
      10'b1001001110 : begin
        result = input_590;
      end
      10'b1001001111 : begin
        result = input_591;
      end
      10'b1001010000 : begin
        result = input_592;
      end
      10'b1001010001 : begin
        result = input_593;
      end
      10'b1001010010 : begin
        result = input_594;
      end
      10'b1001010011 : begin
        result = input_595;
      end
      10'b1001010100 : begin
        result = input_596;
      end
      10'b1001010101 : begin
        result = input_597;
      end
      10'b1001010110 : begin
        result = input_598;
      end
      10'b1001010111 : begin
        result = input_599;
      end
      10'b1001011000 : begin
        result = input_600;
      end
      10'b1001011001 : begin
        result = input_601;
      end
      10'b1001011010 : begin
        result = input_602;
      end
      10'b1001011011 : begin
        result = input_603;
      end
      10'b1001011100 : begin
        result = input_604;
      end
      10'b1001011101 : begin
        result = input_605;
      end
      10'b1001011110 : begin
        result = input_606;
      end
      10'b1001011111 : begin
        result = input_607;
      end
      10'b1001100000 : begin
        result = input_608;
      end
      10'b1001100001 : begin
        result = input_609;
      end
      10'b1001100010 : begin
        result = input_610;
      end
      10'b1001100011 : begin
        result = input_611;
      end
      10'b1001100100 : begin
        result = input_612;
      end
      10'b1001100101 : begin
        result = input_613;
      end
      10'b1001100110 : begin
        result = input_614;
      end
      10'b1001100111 : begin
        result = input_615;
      end
      10'b1001101000 : begin
        result = input_616;
      end
      10'b1001101001 : begin
        result = input_617;
      end
      10'b1001101010 : begin
        result = input_618;
      end
      10'b1001101011 : begin
        result = input_619;
      end
      10'b1001101100 : begin
        result = input_620;
      end
      10'b1001101101 : begin
        result = input_621;
      end
      10'b1001101110 : begin
        result = input_622;
      end
      10'b1001101111 : begin
        result = input_623;
      end
      10'b1001110000 : begin
        result = input_624;
      end
      10'b1001110001 : begin
        result = input_625;
      end
      10'b1001110010 : begin
        result = input_626;
      end
      10'b1001110011 : begin
        result = input_627;
      end
      10'b1001110100 : begin
        result = input_628;
      end
      10'b1001110101 : begin
        result = input_629;
      end
      10'b1001110110 : begin
        result = input_630;
      end
      10'b1001110111 : begin
        result = input_631;
      end
      10'b1001111000 : begin
        result = input_632;
      end
      10'b1001111001 : begin
        result = input_633;
      end
      10'b1001111010 : begin
        result = input_634;
      end
      10'b1001111011 : begin
        result = input_635;
      end
      10'b1001111100 : begin
        result = input_636;
      end
      10'b1001111101 : begin
        result = input_637;
      end
      10'b1001111110 : begin
        result = input_638;
      end
      10'b1001111111 : begin
        result = input_639;
      end
      10'b1010000000 : begin
        result = input_640;
      end
      10'b1010000001 : begin
        result = input_641;
      end
      10'b1010000010 : begin
        result = input_642;
      end
      10'b1010000011 : begin
        result = input_643;
      end
      10'b1010000100 : begin
        result = input_644;
      end
      10'b1010000101 : begin
        result = input_645;
      end
      10'b1010000110 : begin
        result = input_646;
      end
      10'b1010000111 : begin
        result = input_647;
      end
      10'b1010001000 : begin
        result = input_648;
      end
      10'b1010001001 : begin
        result = input_649;
      end
      10'b1010001010 : begin
        result = input_650;
      end
      10'b1010001011 : begin
        result = input_651;
      end
      10'b1010001100 : begin
        result = input_652;
      end
      10'b1010001101 : begin
        result = input_653;
      end
      10'b1010001110 : begin
        result = input_654;
      end
      10'b1010001111 : begin
        result = input_655;
      end
      10'b1010010000 : begin
        result = input_656;
      end
      10'b1010010001 : begin
        result = input_657;
      end
      10'b1010010010 : begin
        result = input_658;
      end
      10'b1010010011 : begin
        result = input_659;
      end
      10'b1010010100 : begin
        result = input_660;
      end
      10'b1010010101 : begin
        result = input_661;
      end
      10'b1010010110 : begin
        result = input_662;
      end
      10'b1010010111 : begin
        result = input_663;
      end
      10'b1010011000 : begin
        result = input_664;
      end
      10'b1010011001 : begin
        result = input_665;
      end
      10'b1010011010 : begin
        result = input_666;
      end
      10'b1010011011 : begin
        result = input_667;
      end
      10'b1010011100 : begin
        result = input_668;
      end
      10'b1010011101 : begin
        result = input_669;
      end
      10'b1010011110 : begin
        result = input_670;
      end
      10'b1010011111 : begin
        result = input_671;
      end
      10'b1010100000 : begin
        result = input_672;
      end
      10'b1010100001 : begin
        result = input_673;
      end
      10'b1010100010 : begin
        result = input_674;
      end
      10'b1010100011 : begin
        result = input_675;
      end
      10'b1010100100 : begin
        result = input_676;
      end
      10'b1010100101 : begin
        result = input_677;
      end
      10'b1010100110 : begin
        result = input_678;
      end
      10'b1010100111 : begin
        result = input_679;
      end
      10'b1010101000 : begin
        result = input_680;
      end
      10'b1010101001 : begin
        result = input_681;
      end
      10'b1010101010 : begin
        result = input_682;
      end
      10'b1010101011 : begin
        result = input_683;
      end
      10'b1010101100 : begin
        result = input_684;
      end
      10'b1010101101 : begin
        result = input_685;
      end
      10'b1010101110 : begin
        result = input_686;
      end
      10'b1010101111 : begin
        result = input_687;
      end
      10'b1010110000 : begin
        result = input_688;
      end
      10'b1010110001 : begin
        result = input_689;
      end
      10'b1010110010 : begin
        result = input_690;
      end
      10'b1010110011 : begin
        result = input_691;
      end
      10'b1010110100 : begin
        result = input_692;
      end
      10'b1010110101 : begin
        result = input_693;
      end
      10'b1010110110 : begin
        result = input_694;
      end
      10'b1010110111 : begin
        result = input_695;
      end
      10'b1010111000 : begin
        result = input_696;
      end
      10'b1010111001 : begin
        result = input_697;
      end
      10'b1010111010 : begin
        result = input_698;
      end
      10'b1010111011 : begin
        result = input_699;
      end
      10'b1010111100 : begin
        result = input_700;
      end
      10'b1010111101 : begin
        result = input_701;
      end
      10'b1010111110 : begin
        result = input_702;
      end
      10'b1010111111 : begin
        result = input_703;
      end
      10'b1011000000 : begin
        result = input_704;
      end
      10'b1011000001 : begin
        result = input_705;
      end
      10'b1011000010 : begin
        result = input_706;
      end
      10'b1011000011 : begin
        result = input_707;
      end
      10'b1011000100 : begin
        result = input_708;
      end
      10'b1011000101 : begin
        result = input_709;
      end
      10'b1011000110 : begin
        result = input_710;
      end
      10'b1011000111 : begin
        result = input_711;
      end
      10'b1011001000 : begin
        result = input_712;
      end
      10'b1011001001 : begin
        result = input_713;
      end
      10'b1011001010 : begin
        result = input_714;
      end
      10'b1011001011 : begin
        result = input_715;
      end
      10'b1011001100 : begin
        result = input_716;
      end
      10'b1011001101 : begin
        result = input_717;
      end
      10'b1011001110 : begin
        result = input_718;
      end
      10'b1011001111 : begin
        result = input_719;
      end
      10'b1011010000 : begin
        result = input_720;
      end
      10'b1011010001 : begin
        result = input_721;
      end
      10'b1011010010 : begin
        result = input_722;
      end
      10'b1011010011 : begin
        result = input_723;
      end
      10'b1011010100 : begin
        result = input_724;
      end
      10'b1011010101 : begin
        result = input_725;
      end
      10'b1011010110 : begin
        result = input_726;
      end
      10'b1011010111 : begin
        result = input_727;
      end
      10'b1011011000 : begin
        result = input_728;
      end
      10'b1011011001 : begin
        result = input_729;
      end
      10'b1011011010 : begin
        result = input_730;
      end
      10'b1011011011 : begin
        result = input_731;
      end
      10'b1011011100 : begin
        result = input_732;
      end
      10'b1011011101 : begin
        result = input_733;
      end
      10'b1011011110 : begin
        result = input_734;
      end
      10'b1011011111 : begin
        result = input_735;
      end
      10'b1011100000 : begin
        result = input_736;
      end
      10'b1011100001 : begin
        result = input_737;
      end
      10'b1011100010 : begin
        result = input_738;
      end
      10'b1011100011 : begin
        result = input_739;
      end
      10'b1011100100 : begin
        result = input_740;
      end
      10'b1011100101 : begin
        result = input_741;
      end
      10'b1011100110 : begin
        result = input_742;
      end
      10'b1011100111 : begin
        result = input_743;
      end
      10'b1011101000 : begin
        result = input_744;
      end
      10'b1011101001 : begin
        result = input_745;
      end
      10'b1011101010 : begin
        result = input_746;
      end
      10'b1011101011 : begin
        result = input_747;
      end
      10'b1011101100 : begin
        result = input_748;
      end
      10'b1011101101 : begin
        result = input_749;
      end
      10'b1011101110 : begin
        result = input_750;
      end
      10'b1011101111 : begin
        result = input_751;
      end
      10'b1011110000 : begin
        result = input_752;
      end
      10'b1011110001 : begin
        result = input_753;
      end
      10'b1011110010 : begin
        result = input_754;
      end
      10'b1011110011 : begin
        result = input_755;
      end
      10'b1011110100 : begin
        result = input_756;
      end
      10'b1011110101 : begin
        result = input_757;
      end
      10'b1011110110 : begin
        result = input_758;
      end
      10'b1011110111 : begin
        result = input_759;
      end
      10'b1011111000 : begin
        result = input_760;
      end
      10'b1011111001 : begin
        result = input_761;
      end
      10'b1011111010 : begin
        result = input_762;
      end
      10'b1011111011 : begin
        result = input_763;
      end
      10'b1011111100 : begin
        result = input_764;
      end
      10'b1011111101 : begin
        result = input_765;
      end
      10'b1011111110 : begin
        result = input_766;
      end
      10'b1011111111 : begin
        result = input_767;
      end
      10'b1100000000 : begin
        result = input_768;
      end
      10'b1100000001 : begin
        result = input_769;
      end
      10'b1100000010 : begin
        result = input_770;
      end
      10'b1100000011 : begin
        result = input_771;
      end
      10'b1100000100 : begin
        result = input_772;
      end
      10'b1100000101 : begin
        result = input_773;
      end
      10'b1100000110 : begin
        result = input_774;
      end
      10'b1100000111 : begin
        result = input_775;
      end
      10'b1100001000 : begin
        result = input_776;
      end
      10'b1100001001 : begin
        result = input_777;
      end
      10'b1100001010 : begin
        result = input_778;
      end
      10'b1100001011 : begin
        result = input_779;
      end
      10'b1100001100 : begin
        result = input_780;
      end
      10'b1100001101 : begin
        result = input_781;
      end
      10'b1100001110 : begin
        result = input_782;
      end
      default : begin
        result = input_783;
      end
    endcase
    MUX_v_18_784_2 = result;
  end
  endfunction


  function automatic [18:0] MUX_v_19_2_2;
    input [18:0] input_0;
    input [18:0] input_1;
    input [0:0] sel;
    reg [18:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_19_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_64_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [1:0] input_2;
    input [1:0] input_3;
    input [1:0] input_4;
    input [1:0] input_5;
    input [1:0] input_6;
    input [1:0] input_7;
    input [1:0] input_8;
    input [1:0] input_9;
    input [1:0] input_10;
    input [1:0] input_11;
    input [1:0] input_12;
    input [1:0] input_13;
    input [1:0] input_14;
    input [1:0] input_15;
    input [1:0] input_16;
    input [1:0] input_17;
    input [1:0] input_18;
    input [1:0] input_19;
    input [1:0] input_20;
    input [1:0] input_21;
    input [1:0] input_22;
    input [1:0] input_23;
    input [1:0] input_24;
    input [1:0] input_25;
    input [1:0] input_26;
    input [1:0] input_27;
    input [1:0] input_28;
    input [1:0] input_29;
    input [1:0] input_30;
    input [1:0] input_31;
    input [1:0] input_32;
    input [1:0] input_33;
    input [1:0] input_34;
    input [1:0] input_35;
    input [1:0] input_36;
    input [1:0] input_37;
    input [1:0] input_38;
    input [1:0] input_39;
    input [1:0] input_40;
    input [1:0] input_41;
    input [1:0] input_42;
    input [1:0] input_43;
    input [1:0] input_44;
    input [1:0] input_45;
    input [1:0] input_46;
    input [1:0] input_47;
    input [1:0] input_48;
    input [1:0] input_49;
    input [1:0] input_50;
    input [1:0] input_51;
    input [1:0] input_52;
    input [1:0] input_53;
    input [1:0] input_54;
    input [1:0] input_55;
    input [1:0] input_56;
    input [1:0] input_57;
    input [1:0] input_58;
    input [1:0] input_59;
    input [1:0] input_60;
    input [1:0] input_61;
    input [1:0] input_62;
    input [1:0] input_63;
    input [5:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_2_64_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_4_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [2:0] input_2;
    input [2:0] input_3;
    input [1:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_3_4_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_4_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [4:0] input_2;
    input [4:0] input_3;
    input [1:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_5_4_2 = result;
  end
  endfunction


  function automatic [67:0] MUX_v_68_2_2;
    input [67:0] input_0;
    input [67:0] input_1;
    input [0:0] sel;
    reg [67:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_68_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_16_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [5:0] input_2;
    input [5:0] input_3;
    input [5:0] input_4;
    input [5:0] input_5;
    input [5:0] input_6;
    input [5:0] input_7;
    input [5:0] input_8;
    input [5:0] input_9;
    input [5:0] input_10;
    input [5:0] input_11;
    input [5:0] input_12;
    input [5:0] input_13;
    input [5:0] input_14;
    input [5:0] input_15;
    input [3:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_6_16_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [69:0] MUX_v_70_2_2;
    input [69:0] input_0;
    input [69:0] input_1;
    input [0:0] sel;
    reg [69:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_70_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_4_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [6:0] input_2;
    input [6:0] input_3;
    input [1:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_7_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [90:0] MUX_v_91_2_2;
    input [90:0] input_0;
    input [90:0] input_1;
    input [0:0] sel;
    reg [90:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_91_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [147:0] readslicef_158_148_10;
    input [157:0] vector;
    reg [157:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_158_148_10 = tmp[147:0];
  end
  endfunction


  function automatic [14:0] readslicef_23_15_8;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_23_15_8 = tmp[14:0];
  end
  endfunction


  function automatic [17:0] readslicef_28_18_10;
    input [27:0] vector;
    reg [27:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_28_18_10 = tmp[17:0];
  end
  endfunction


  function automatic [0:0] readslicef_4_1_3;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_4_1_3 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_7_1_6;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_7_1_6 = tmp[0:0];
  end
  endfunction


  function automatic [6:0] readslicef_8_7_1;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_8_7_1 = tmp[6:0];
  end
  endfunction


  function automatic [9:0] signext_10_1;
    input [0:0] vector;
  begin
    signext_10_1= {{9{vector[0]}}, vector};
  end
  endfunction


  function automatic [14:0] signext_15_10;
    input [9:0] vector;
  begin
    signext_15_10= {{5{vector[9]}}, vector};
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input [0:0] vector;
  begin
    signext_2_1= {{1{vector[0]}}, vector};
  end
  endfunction


  function automatic [2:0] signext_3_1;
    input [0:0] vector;
  begin
    signext_3_1= {{2{vector[0]}}, vector};
  end
  endfunction


  function automatic [3:0] signext_4_1;
    input [0:0] vector;
  begin
    signext_4_1= {{3{vector[0]}}, vector};
  end
  endfunction


  function automatic [73:0] signext_74_1;
    input [0:0] vector;
  begin
    signext_74_1= {{73{vector[0]}}, vector};
  end
  endfunction


  function automatic [7:0] signext_8_4;
    input [3:0] vector;
  begin
    signext_8_4= {{4{vector[3]}}, vector};
  end
  endfunction


  function automatic [5:0] conv_s2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_s2u_5_6 = {vector[4], vector};
  end
  endfunction


  function automatic [8:0] conv_s2u_7_9 ;
    input [6:0]  vector ;
  begin
    conv_s2u_7_9 = {{2{vector[6]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_s2u_9_11 ;
    input [8:0]  vector ;
  begin
    conv_s2u_9_11 = {{2{vector[8]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_15_18 ;
    input [14:0]  vector ;
  begin
    conv_s2u_15_18 = {{3{vector[14]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_16_19 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_19 = {{3{vector[15]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_17_19 ;
    input [16:0]  vector ;
  begin
    conv_s2u_17_19 = {{2{vector[16]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_19 = {vector[17], vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_18_22 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_22 = {{4{vector[17]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2u_19_20 ;
    input [18:0]  vector ;
  begin
    conv_s2u_19_20 = {vector[18], vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_21_22 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_22 = {vector[20], vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_21_23 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_23 = {{2{vector[20]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_22_23 ;
    input [21:0]  vector ;
  begin
    conv_s2u_22_23 = {vector[21], vector};
  end
  endfunction


  function automatic [5:0] conv_u2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2s_5_6 =  {1'b0, vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_7 =  {1'b0, vector};
  end
  endfunction


  function automatic [17:0] conv_u2s_17_18 ;
    input [16:0]  vector ;
  begin
    conv_u2s_17_18 =  {1'b0, vector};
  end
  endfunction


  function automatic [67:0] conv_u2s_67_68 ;
    input [66:0]  vector ;
  begin
    conv_u2s_67_68 =  {1'b0, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_1_4 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_4 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_1_8 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_8 = {{7{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_2_8 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_8 = {{6{1'b0}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_5_7 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_7 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_5_8 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_8 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_6_8 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_8 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_9_11 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_11 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [18:0] conv_u2u_19_19 ;
    input [18:0]  vector ;
  begin
    conv_u2u_19_19 = vector;
  end
  endfunction


  function automatic [67:0] conv_u2u_67_68 ;
    input [66:0]  vector ;
  begin
    conv_u2u_67_68 = {1'b0, vector};
  end
  endfunction


  function automatic [68:0] conv_u2u_68_69 ;
    input [67:0]  vector ;
  begin
    conv_u2u_68_69 = {1'b0, vector};
  end
  endfunction


  function automatic [70:0] conv_u2u_69_71 ;
    input [68:0]  vector ;
  begin
    conv_u2u_69_71 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [70:0] conv_u2u_70_71 ;
    input [69:0]  vector ;
  begin
    conv_u2u_70_71 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    mnist_mlp
// ------------------------------------------------------------------


module mnist_mlp (
  clk, rst, 
  
  // Input Feature
  input1_rsc_dat, input1_rsc_vld, input1_rsc_rdy,
  
  // Prediction
  layer7_out_rsc_dat, layer7_out_rsc_vld, layer7_out_rsc_rdy,
  
  // Some I/O constants (ignore)
  const_size_in_1_rsc_dat, const_size_in_1_rsc_vld, const_size_in_1_rsc_rdy,
  const_size_out_1_rsc_dat, const_size_out_1_rsc_vld, const_size_out_1_rsc_rdy,

  // Weights and biases in external SRAMs
  w2_rsc_adra, w2_rsc_da, w2_rsc_ena, w2_rsc_wea, w2_rsc_qa, w2_rsc_adrb, w2_rsc_db, w2_rsc_enb, w2_rsc_web, w2_rsc_qb,
  b2_rsc_dat,
  w4_rsc_adra, w4_rsc_da, w4_rsc_ena, w4_rsc_wea, w4_rsc_qa, w4_rsc_adrb, w4_rsc_db, w4_rsc_enb, w4_rsc_web, w4_rsc_qb,
  b4_rsc_dat,
  w6_rsc_adra, w6_rsc_da, w6_rsc_ena, w6_rsc_wea, w6_rsc_qa, w6_rsc_adrb, w6_rsc_db, w6_rsc_enb, w6_rsc_web, w6_rsc_qb,
  b6_rsc_dat
);
  input clk;
  input rst;
  input [14111:0] input1_rsc_dat;
  input input1_rsc_vld;
  output input1_rsc_rdy;
  output [179:0] layer7_out_rsc_dat;
  output layer7_out_rsc_vld;
  input layer7_out_rsc_rdy;
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  input const_size_in_1_rsc_rdy;
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  input const_size_out_1_rsc_rdy;
  output [15:0] w2_rsc_adra;
  output [17:0] w2_rsc_da;
  output w2_rsc_ena;
  output w2_rsc_wea;
  input [17:0] w2_rsc_qa;
  output [15:0] w2_rsc_adrb;
  output [17:0] w2_rsc_db;
  output w2_rsc_enb;
  output w2_rsc_web;
  input [17:0] w2_rsc_qb;
  input [1151:0] b2_rsc_dat;
  output [11:0] w4_rsc_adra;
  output [17:0] w4_rsc_da;
  output w4_rsc_ena;
  output w4_rsc_wea;
  input [17:0] w4_rsc_qa;
  output [11:0] w4_rsc_adrb;
  output [17:0] w4_rsc_db;
  output w4_rsc_enb;
  output w4_rsc_web;
  input [17:0] w4_rsc_qb;
  input [1151:0] b4_rsc_dat;
  output [9:0] w6_rsc_adra;
  output [17:0] w6_rsc_da;
  output w6_rsc_ena;
  output w6_rsc_wea;
  input [17:0] w6_rsc_qa;
  output [9:0] w6_rsc_adrb;
  output [17:0] w6_rsc_db;
  output w6_rsc_enb;
  output w6_rsc_web;
  input [17:0] w6_rsc_qb;
  input [179:0] b6_rsc_dat;


  // Interconnect Declarations
  wire [31:0] w2_rsci_adra_d;
  wire [1:0] w2_rsci_ena_d;
  wire [35:0] w2_rsci_qa_d;
  wire [1:0] w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [23:0] w4_rsci_adra_d;
  wire [1:0] w4_rsci_ena_d;
  wire [35:0] w4_rsci_qa_d;
  wire [1:0] w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [19:0] w6_rsci_adra_d;
  wire [1:0] w6_rsci_ena_d;
  wire [35:0] w6_rsci_qa_d;
  wire [1:0] w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations for Component Instantiations 
  mnist_mlp_ccs_sample_mem_ccs_ram_sync_dualport_rwport_5_18_16_50176_50176_18_5_gen
      w2_rsci (
      .qb(w2_rsc_qb),
      .web(w2_rsc_web),
      .enb(w2_rsc_enb),
      .db(w2_rsc_db),
      .adrb(w2_rsc_adrb),
      .qa(w2_rsc_qa),
      .wea(w2_rsc_wea),
      .ena(w2_rsc_ena),
      .da(w2_rsc_da),
      .adra(w2_rsc_adra),
      .adra_d(w2_rsci_adra_d),
      .da_d(36'b000000000000000000000000000000000000),
      .ena_d(w2_rsci_ena_d),
      .wea_d(2'b00),
      .qa_d(w2_rsci_qa_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  mnist_mlp_ccs_sample_mem_ccs_ram_sync_dualport_rwport_7_18_12_4096_4096_18_5_gen
      w4_rsci (
      .qb(w4_rsc_qb),
      .web(w4_rsc_web),
      .enb(w4_rsc_enb),
      .db(w4_rsc_db),
      .adrb(w4_rsc_adrb),
      .qa(w4_rsc_qa),
      .wea(w4_rsc_wea),
      .ena(w4_rsc_ena),
      .da(w4_rsc_da),
      .adra(w4_rsc_adra),
      .adra_d(w4_rsci_adra_d),
      .da_d(36'b000000000000000000000000000000000000),
      .ena_d(w4_rsci_ena_d),
      .wea_d(2'b00),
      .qa_d(w4_rsci_qa_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  mnist_mlp_ccs_sample_mem_ccs_ram_sync_dualport_rwport_9_18_10_640_640_18_5_gen
      w6_rsci (
      .qb(w6_rsc_qb),
      .web(w6_rsc_web),
      .enb(w6_rsc_enb),
      .db(w6_rsc_db),
      .adrb(w6_rsc_adrb),
      .qa(w6_rsc_qa),
      .wea(w6_rsc_wea),
      .ena(w6_rsc_ena),
      .da(w6_rsc_da),
      .adra(w6_rsc_adra),
      .adra_d(w6_rsci_adra_d),
      .da_d(36'b000000000000000000000000000000000000),
      .ena_d(w6_rsci_ena_d),
      .wea_d(2'b00),
      .qa_d(w6_rsci_qa_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  mnist_mlp_core mnist_mlp_core_inst (
      .clk(clk),
      .rst(rst),
      .input1_rsc_dat(input1_rsc_dat),
      .input1_rsc_vld(input1_rsc_vld),
      .input1_rsc_rdy(input1_rsc_rdy),
      .layer7_out_rsc_dat(layer7_out_rsc_dat),
      .layer7_out_rsc_vld(layer7_out_rsc_vld),
      .layer7_out_rsc_rdy(layer7_out_rsc_rdy),
      .const_size_in_1_rsc_dat(const_size_in_1_rsc_dat),
      .const_size_in_1_rsc_vld(const_size_in_1_rsc_vld),
      .const_size_in_1_rsc_rdy(const_size_in_1_rsc_rdy),
      .const_size_out_1_rsc_dat(const_size_out_1_rsc_dat),
      .const_size_out_1_rsc_vld(const_size_out_1_rsc_vld),
      .const_size_out_1_rsc_rdy(const_size_out_1_rsc_rdy),
      .b2_rsc_dat(b2_rsc_dat),
      .b4_rsc_dat(b4_rsc_dat),
      .b6_rsc_dat(b6_rsc_dat),
      .w2_rsci_adra_d(w2_rsci_adra_d),
      .w2_rsci_ena_d(w2_rsci_ena_d),
      .w2_rsci_qa_d(w2_rsci_qa_d),
      .w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(w2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .w4_rsci_adra_d(w4_rsci_adra_d),
      .w4_rsci_ena_d(w4_rsci_ena_d),
      .w4_rsci_qa_d(w4_rsci_qa_d),
      .w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(w4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .w6_rsci_adra_d(w6_rsci_adra_d),
      .w6_rsci_ena_d(w6_rsci_ena_d),
      .w6_rsci_qa_d(w6_rsci_qa_d),
      .w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(w6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d)
    );
endmodule



