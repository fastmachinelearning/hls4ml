//----------------------------------------------------------------------
//----------------------------------------------------------------------
// Created by      : giuseppe
// Creation Date   : 2019 Dec 05
// Created with uvmf_gen version 2019.1
//----------------------------------------------------------------------
//
//----------------------------------------------------------------------
// Project         : mnist_mlp_bench Simulation Bench 
// Unit            : Top level UVM test
// File            : test_top.svh
//----------------------------------------------------------------------
// Description: This top level UVM test is the base class for all
//     future tests created for this project.
//
//     This test class contains:
//          Configuration:  The top level configuration for the project.
//          Environment:    The top level environment for the project.
//          Top_level_sequence:  The top level sequence for the project.
//                                       f   
//----------------------------------------------------------------------
//

typedef mnist_mlp_env_configuration mnist_mlp_env_configuration_t;
typedef mnist_mlp_environment mnist_mlp_environment_t;

class test_top extends uvmf_test_base #(.CONFIG_T(mnist_mlp_env_configuration_t), 
                                        .ENV_T(mnist_mlp_environment_t), 
                                        .TOP_LEVEL_SEQ_T(mnist_mlp_bench_bench_sequence_base));

  `uvm_component_utils( test_top );


  string interface_names[] = {
    input1_rsc_BFM /* input1_rsc     [0] */ , 
    output1_rsc_BFM /* output1_rsc     [1] */ , 
    const_size_in_1_rsc_BFM /* const_size_in_1_rsc     [2] */ , 
    const_size_out_1_rsc_BFM /* const_size_out_1_rsc     [3] */ , 
    w2_rsc_0_0_BFM /* w2_rsc_0_0     [4] */ , 
    w2_rsc_1_0_BFM /* w2_rsc_1_0     [5] */ , 
    w2_rsc_2_0_BFM /* w2_rsc_2_0     [6] */ , 
    w2_rsc_3_0_BFM /* w2_rsc_3_0     [7] */ , 
    w2_rsc_4_0_BFM /* w2_rsc_4_0     [8] */ , 
    w2_rsc_5_0_BFM /* w2_rsc_5_0     [9] */ , 
    w2_rsc_6_0_BFM /* w2_rsc_6_0     [10] */ , 
    w2_rsc_7_0_BFM /* w2_rsc_7_0     [11] */ , 
    w2_rsc_8_0_BFM /* w2_rsc_8_0     [12] */ , 
    w2_rsc_9_0_BFM /* w2_rsc_9_0     [13] */ , 
    w2_rsc_10_0_BFM /* w2_rsc_10_0     [14] */ , 
    w2_rsc_11_0_BFM /* w2_rsc_11_0     [15] */ , 
    w2_rsc_12_0_BFM /* w2_rsc_12_0     [16] */ , 
    w2_rsc_13_0_BFM /* w2_rsc_13_0     [17] */ , 
    w2_rsc_14_0_BFM /* w2_rsc_14_0     [18] */ , 
    w2_rsc_15_0_BFM /* w2_rsc_15_0     [19] */ , 
    w2_rsc_16_0_BFM /* w2_rsc_16_0     [20] */ , 
    w2_rsc_17_0_BFM /* w2_rsc_17_0     [21] */ , 
    w2_rsc_18_0_BFM /* w2_rsc_18_0     [22] */ , 
    w2_rsc_19_0_BFM /* w2_rsc_19_0     [23] */ , 
    w2_rsc_20_0_BFM /* w2_rsc_20_0     [24] */ , 
    w2_rsc_21_0_BFM /* w2_rsc_21_0     [25] */ , 
    w2_rsc_22_0_BFM /* w2_rsc_22_0     [26] */ , 
    w2_rsc_23_0_BFM /* w2_rsc_23_0     [27] */ , 
    w2_rsc_24_0_BFM /* w2_rsc_24_0     [28] */ , 
    w2_rsc_25_0_BFM /* w2_rsc_25_0     [29] */ , 
    w2_rsc_26_0_BFM /* w2_rsc_26_0     [30] */ , 
    w2_rsc_27_0_BFM /* w2_rsc_27_0     [31] */ , 
    w2_rsc_28_0_BFM /* w2_rsc_28_0     [32] */ , 
    w2_rsc_29_0_BFM /* w2_rsc_29_0     [33] */ , 
    w2_rsc_30_0_BFM /* w2_rsc_30_0     [34] */ , 
    w2_rsc_31_0_BFM /* w2_rsc_31_0     [35] */ , 
    w2_rsc_32_0_BFM /* w2_rsc_32_0     [36] */ , 
    w2_rsc_33_0_BFM /* w2_rsc_33_0     [37] */ , 
    w2_rsc_34_0_BFM /* w2_rsc_34_0     [38] */ , 
    w2_rsc_35_0_BFM /* w2_rsc_35_0     [39] */ , 
    w2_rsc_36_0_BFM /* w2_rsc_36_0     [40] */ , 
    w2_rsc_37_0_BFM /* w2_rsc_37_0     [41] */ , 
    w2_rsc_38_0_BFM /* w2_rsc_38_0     [42] */ , 
    w2_rsc_39_0_BFM /* w2_rsc_39_0     [43] */ , 
    w2_rsc_40_0_BFM /* w2_rsc_40_0     [44] */ , 
    w2_rsc_41_0_BFM /* w2_rsc_41_0     [45] */ , 
    w2_rsc_42_0_BFM /* w2_rsc_42_0     [46] */ , 
    w2_rsc_43_0_BFM /* w2_rsc_43_0     [47] */ , 
    w2_rsc_44_0_BFM /* w2_rsc_44_0     [48] */ , 
    w2_rsc_45_0_BFM /* w2_rsc_45_0     [49] */ , 
    w2_rsc_46_0_BFM /* w2_rsc_46_0     [50] */ , 
    w2_rsc_47_0_BFM /* w2_rsc_47_0     [51] */ , 
    w2_rsc_48_0_BFM /* w2_rsc_48_0     [52] */ , 
    w2_rsc_49_0_BFM /* w2_rsc_49_0     [53] */ , 
    w2_rsc_50_0_BFM /* w2_rsc_50_0     [54] */ , 
    w2_rsc_51_0_BFM /* w2_rsc_51_0     [55] */ , 
    w2_rsc_52_0_BFM /* w2_rsc_52_0     [56] */ , 
    w2_rsc_53_0_BFM /* w2_rsc_53_0     [57] */ , 
    w2_rsc_54_0_BFM /* w2_rsc_54_0     [58] */ , 
    w2_rsc_55_0_BFM /* w2_rsc_55_0     [59] */ , 
    w2_rsc_56_0_BFM /* w2_rsc_56_0     [60] */ , 
    w2_rsc_57_0_BFM /* w2_rsc_57_0     [61] */ , 
    w2_rsc_58_0_BFM /* w2_rsc_58_0     [62] */ , 
    w2_rsc_59_0_BFM /* w2_rsc_59_0     [63] */ , 
    w2_rsc_60_0_BFM /* w2_rsc_60_0     [64] */ , 
    w2_rsc_61_0_BFM /* w2_rsc_61_0     [65] */ , 
    w2_rsc_62_0_BFM /* w2_rsc_62_0     [66] */ , 
    w2_rsc_63_0_BFM /* w2_rsc_63_0     [67] */ , 
    b2_rsc_BFM /* b2_rsc     [68] */ , 
    w4_rsc_0_0_BFM /* w4_rsc_0_0     [69] */ , 
    w4_rsc_1_0_BFM /* w4_rsc_1_0     [70] */ , 
    w4_rsc_2_0_BFM /* w4_rsc_2_0     [71] */ , 
    w4_rsc_3_0_BFM /* w4_rsc_3_0     [72] */ , 
    w4_rsc_4_0_BFM /* w4_rsc_4_0     [73] */ , 
    w4_rsc_5_0_BFM /* w4_rsc_5_0     [74] */ , 
    w4_rsc_6_0_BFM /* w4_rsc_6_0     [75] */ , 
    w4_rsc_7_0_BFM /* w4_rsc_7_0     [76] */ , 
    w4_rsc_8_0_BFM /* w4_rsc_8_0     [77] */ , 
    w4_rsc_9_0_BFM /* w4_rsc_9_0     [78] */ , 
    w4_rsc_10_0_BFM /* w4_rsc_10_0     [79] */ , 
    w4_rsc_11_0_BFM /* w4_rsc_11_0     [80] */ , 
    w4_rsc_12_0_BFM /* w4_rsc_12_0     [81] */ , 
    w4_rsc_13_0_BFM /* w4_rsc_13_0     [82] */ , 
    w4_rsc_14_0_BFM /* w4_rsc_14_0     [83] */ , 
    w4_rsc_15_0_BFM /* w4_rsc_15_0     [84] */ , 
    w4_rsc_16_0_BFM /* w4_rsc_16_0     [85] */ , 
    w4_rsc_17_0_BFM /* w4_rsc_17_0     [86] */ , 
    w4_rsc_18_0_BFM /* w4_rsc_18_0     [87] */ , 
    w4_rsc_19_0_BFM /* w4_rsc_19_0     [88] */ , 
    w4_rsc_20_0_BFM /* w4_rsc_20_0     [89] */ , 
    w4_rsc_21_0_BFM /* w4_rsc_21_0     [90] */ , 
    w4_rsc_22_0_BFM /* w4_rsc_22_0     [91] */ , 
    w4_rsc_23_0_BFM /* w4_rsc_23_0     [92] */ , 
    w4_rsc_24_0_BFM /* w4_rsc_24_0     [93] */ , 
    w4_rsc_25_0_BFM /* w4_rsc_25_0     [94] */ , 
    w4_rsc_26_0_BFM /* w4_rsc_26_0     [95] */ , 
    w4_rsc_27_0_BFM /* w4_rsc_27_0     [96] */ , 
    w4_rsc_28_0_BFM /* w4_rsc_28_0     [97] */ , 
    w4_rsc_29_0_BFM /* w4_rsc_29_0     [98] */ , 
    w4_rsc_30_0_BFM /* w4_rsc_30_0     [99] */ , 
    w4_rsc_31_0_BFM /* w4_rsc_31_0     [100] */ , 
    w4_rsc_32_0_BFM /* w4_rsc_32_0     [101] */ , 
    w4_rsc_33_0_BFM /* w4_rsc_33_0     [102] */ , 
    w4_rsc_34_0_BFM /* w4_rsc_34_0     [103] */ , 
    w4_rsc_35_0_BFM /* w4_rsc_35_0     [104] */ , 
    w4_rsc_36_0_BFM /* w4_rsc_36_0     [105] */ , 
    w4_rsc_37_0_BFM /* w4_rsc_37_0     [106] */ , 
    w4_rsc_38_0_BFM /* w4_rsc_38_0     [107] */ , 
    w4_rsc_39_0_BFM /* w4_rsc_39_0     [108] */ , 
    w4_rsc_40_0_BFM /* w4_rsc_40_0     [109] */ , 
    w4_rsc_41_0_BFM /* w4_rsc_41_0     [110] */ , 
    w4_rsc_42_0_BFM /* w4_rsc_42_0     [111] */ , 
    w4_rsc_43_0_BFM /* w4_rsc_43_0     [112] */ , 
    w4_rsc_44_0_BFM /* w4_rsc_44_0     [113] */ , 
    w4_rsc_45_0_BFM /* w4_rsc_45_0     [114] */ , 
    w4_rsc_46_0_BFM /* w4_rsc_46_0     [115] */ , 
    w4_rsc_47_0_BFM /* w4_rsc_47_0     [116] */ , 
    w4_rsc_48_0_BFM /* w4_rsc_48_0     [117] */ , 
    w4_rsc_49_0_BFM /* w4_rsc_49_0     [118] */ , 
    w4_rsc_50_0_BFM /* w4_rsc_50_0     [119] */ , 
    w4_rsc_51_0_BFM /* w4_rsc_51_0     [120] */ , 
    w4_rsc_52_0_BFM /* w4_rsc_52_0     [121] */ , 
    w4_rsc_53_0_BFM /* w4_rsc_53_0     [122] */ , 
    w4_rsc_54_0_BFM /* w4_rsc_54_0     [123] */ , 
    w4_rsc_55_0_BFM /* w4_rsc_55_0     [124] */ , 
    w4_rsc_56_0_BFM /* w4_rsc_56_0     [125] */ , 
    w4_rsc_57_0_BFM /* w4_rsc_57_0     [126] */ , 
    w4_rsc_58_0_BFM /* w4_rsc_58_0     [127] */ , 
    w4_rsc_59_0_BFM /* w4_rsc_59_0     [128] */ , 
    w4_rsc_60_0_BFM /* w4_rsc_60_0     [129] */ , 
    w4_rsc_61_0_BFM /* w4_rsc_61_0     [130] */ , 
    w4_rsc_62_0_BFM /* w4_rsc_62_0     [131] */ , 
    w4_rsc_63_0_BFM /* w4_rsc_63_0     [132] */ , 
    b4_rsc_BFM /* b4_rsc     [133] */ , 
    w6_rsc_0_0_BFM /* w6_rsc_0_0     [134] */ , 
    w6_rsc_1_0_BFM /* w6_rsc_1_0     [135] */ , 
    w6_rsc_2_0_BFM /* w6_rsc_2_0     [136] */ , 
    w6_rsc_3_0_BFM /* w6_rsc_3_0     [137] */ , 
    w6_rsc_4_0_BFM /* w6_rsc_4_0     [138] */ , 
    w6_rsc_5_0_BFM /* w6_rsc_5_0     [139] */ , 
    w6_rsc_6_0_BFM /* w6_rsc_6_0     [140] */ , 
    w6_rsc_7_0_BFM /* w6_rsc_7_0     [141] */ , 
    w6_rsc_8_0_BFM /* w6_rsc_8_0     [142] */ , 
    w6_rsc_9_0_BFM /* w6_rsc_9_0     [143] */ , 
    b6_rsc_BFM /* b6_rsc     [144] */ 
};

uvmf_active_passive_t interface_activities[] = { 
    ACTIVE /* input1_rsc     [0] */ , 
    ACTIVE /* output1_rsc     [1] */ , 
    ACTIVE /* const_size_in_1_rsc     [2] */ , 
    ACTIVE /* const_size_out_1_rsc     [3] */ , 
    ACTIVE /* w2_rsc_0_0     [4] */ , 
    ACTIVE /* w2_rsc_1_0     [5] */ , 
    ACTIVE /* w2_rsc_2_0     [6] */ , 
    ACTIVE /* w2_rsc_3_0     [7] */ , 
    ACTIVE /* w2_rsc_4_0     [8] */ , 
    ACTIVE /* w2_rsc_5_0     [9] */ , 
    ACTIVE /* w2_rsc_6_0     [10] */ , 
    ACTIVE /* w2_rsc_7_0     [11] */ , 
    ACTIVE /* w2_rsc_8_0     [12] */ , 
    ACTIVE /* w2_rsc_9_0     [13] */ , 
    ACTIVE /* w2_rsc_10_0     [14] */ , 
    ACTIVE /* w2_rsc_11_0     [15] */ , 
    ACTIVE /* w2_rsc_12_0     [16] */ , 
    ACTIVE /* w2_rsc_13_0     [17] */ , 
    ACTIVE /* w2_rsc_14_0     [18] */ , 
    ACTIVE /* w2_rsc_15_0     [19] */ , 
    ACTIVE /* w2_rsc_16_0     [20] */ , 
    ACTIVE /* w2_rsc_17_0     [21] */ , 
    ACTIVE /* w2_rsc_18_0     [22] */ , 
    ACTIVE /* w2_rsc_19_0     [23] */ , 
    ACTIVE /* w2_rsc_20_0     [24] */ , 
    ACTIVE /* w2_rsc_21_0     [25] */ , 
    ACTIVE /* w2_rsc_22_0     [26] */ , 
    ACTIVE /* w2_rsc_23_0     [27] */ , 
    ACTIVE /* w2_rsc_24_0     [28] */ , 
    ACTIVE /* w2_rsc_25_0     [29] */ , 
    ACTIVE /* w2_rsc_26_0     [30] */ , 
    ACTIVE /* w2_rsc_27_0     [31] */ , 
    ACTIVE /* w2_rsc_28_0     [32] */ , 
    ACTIVE /* w2_rsc_29_0     [33] */ , 
    ACTIVE /* w2_rsc_30_0     [34] */ , 
    ACTIVE /* w2_rsc_31_0     [35] */ , 
    ACTIVE /* w2_rsc_32_0     [36] */ , 
    ACTIVE /* w2_rsc_33_0     [37] */ , 
    ACTIVE /* w2_rsc_34_0     [38] */ , 
    ACTIVE /* w2_rsc_35_0     [39] */ , 
    ACTIVE /* w2_rsc_36_0     [40] */ , 
    ACTIVE /* w2_rsc_37_0     [41] */ , 
    ACTIVE /* w2_rsc_38_0     [42] */ , 
    ACTIVE /* w2_rsc_39_0     [43] */ , 
    ACTIVE /* w2_rsc_40_0     [44] */ , 
    ACTIVE /* w2_rsc_41_0     [45] */ , 
    ACTIVE /* w2_rsc_42_0     [46] */ , 
    ACTIVE /* w2_rsc_43_0     [47] */ , 
    ACTIVE /* w2_rsc_44_0     [48] */ , 
    ACTIVE /* w2_rsc_45_0     [49] */ , 
    ACTIVE /* w2_rsc_46_0     [50] */ , 
    ACTIVE /* w2_rsc_47_0     [51] */ , 
    ACTIVE /* w2_rsc_48_0     [52] */ , 
    ACTIVE /* w2_rsc_49_0     [53] */ , 
    ACTIVE /* w2_rsc_50_0     [54] */ , 
    ACTIVE /* w2_rsc_51_0     [55] */ , 
    ACTIVE /* w2_rsc_52_0     [56] */ , 
    ACTIVE /* w2_rsc_53_0     [57] */ , 
    ACTIVE /* w2_rsc_54_0     [58] */ , 
    ACTIVE /* w2_rsc_55_0     [59] */ , 
    ACTIVE /* w2_rsc_56_0     [60] */ , 
    ACTIVE /* w2_rsc_57_0     [61] */ , 
    ACTIVE /* w2_rsc_58_0     [62] */ , 
    ACTIVE /* w2_rsc_59_0     [63] */ , 
    ACTIVE /* w2_rsc_60_0     [64] */ , 
    ACTIVE /* w2_rsc_61_0     [65] */ , 
    ACTIVE /* w2_rsc_62_0     [66] */ , 
    ACTIVE /* w2_rsc_63_0     [67] */ , 
    ACTIVE /* b2_rsc     [68] */ , 
    ACTIVE /* w4_rsc_0_0     [69] */ , 
    ACTIVE /* w4_rsc_1_0     [70] */ , 
    ACTIVE /* w4_rsc_2_0     [71] */ , 
    ACTIVE /* w4_rsc_3_0     [72] */ , 
    ACTIVE /* w4_rsc_4_0     [73] */ , 
    ACTIVE /* w4_rsc_5_0     [74] */ , 
    ACTIVE /* w4_rsc_6_0     [75] */ , 
    ACTIVE /* w4_rsc_7_0     [76] */ , 
    ACTIVE /* w4_rsc_8_0     [77] */ , 
    ACTIVE /* w4_rsc_9_0     [78] */ , 
    ACTIVE /* w4_rsc_10_0     [79] */ , 
    ACTIVE /* w4_rsc_11_0     [80] */ , 
    ACTIVE /* w4_rsc_12_0     [81] */ , 
    ACTIVE /* w4_rsc_13_0     [82] */ , 
    ACTIVE /* w4_rsc_14_0     [83] */ , 
    ACTIVE /* w4_rsc_15_0     [84] */ , 
    ACTIVE /* w4_rsc_16_0     [85] */ , 
    ACTIVE /* w4_rsc_17_0     [86] */ , 
    ACTIVE /* w4_rsc_18_0     [87] */ , 
    ACTIVE /* w4_rsc_19_0     [88] */ , 
    ACTIVE /* w4_rsc_20_0     [89] */ , 
    ACTIVE /* w4_rsc_21_0     [90] */ , 
    ACTIVE /* w4_rsc_22_0     [91] */ , 
    ACTIVE /* w4_rsc_23_0     [92] */ , 
    ACTIVE /* w4_rsc_24_0     [93] */ , 
    ACTIVE /* w4_rsc_25_0     [94] */ , 
    ACTIVE /* w4_rsc_26_0     [95] */ , 
    ACTIVE /* w4_rsc_27_0     [96] */ , 
    ACTIVE /* w4_rsc_28_0     [97] */ , 
    ACTIVE /* w4_rsc_29_0     [98] */ , 
    ACTIVE /* w4_rsc_30_0     [99] */ , 
    ACTIVE /* w4_rsc_31_0     [100] */ , 
    ACTIVE /* w4_rsc_32_0     [101] */ , 
    ACTIVE /* w4_rsc_33_0     [102] */ , 
    ACTIVE /* w4_rsc_34_0     [103] */ , 
    ACTIVE /* w4_rsc_35_0     [104] */ , 
    ACTIVE /* w4_rsc_36_0     [105] */ , 
    ACTIVE /* w4_rsc_37_0     [106] */ , 
    ACTIVE /* w4_rsc_38_0     [107] */ , 
    ACTIVE /* w4_rsc_39_0     [108] */ , 
    ACTIVE /* w4_rsc_40_0     [109] */ , 
    ACTIVE /* w4_rsc_41_0     [110] */ , 
    ACTIVE /* w4_rsc_42_0     [111] */ , 
    ACTIVE /* w4_rsc_43_0     [112] */ , 
    ACTIVE /* w4_rsc_44_0     [113] */ , 
    ACTIVE /* w4_rsc_45_0     [114] */ , 
    ACTIVE /* w4_rsc_46_0     [115] */ , 
    ACTIVE /* w4_rsc_47_0     [116] */ , 
    ACTIVE /* w4_rsc_48_0     [117] */ , 
    ACTIVE /* w4_rsc_49_0     [118] */ , 
    ACTIVE /* w4_rsc_50_0     [119] */ , 
    ACTIVE /* w4_rsc_51_0     [120] */ , 
    ACTIVE /* w4_rsc_52_0     [121] */ , 
    ACTIVE /* w4_rsc_53_0     [122] */ , 
    ACTIVE /* w4_rsc_54_0     [123] */ , 
    ACTIVE /* w4_rsc_55_0     [124] */ , 
    ACTIVE /* w4_rsc_56_0     [125] */ , 
    ACTIVE /* w4_rsc_57_0     [126] */ , 
    ACTIVE /* w4_rsc_58_0     [127] */ , 
    ACTIVE /* w4_rsc_59_0     [128] */ , 
    ACTIVE /* w4_rsc_60_0     [129] */ , 
    ACTIVE /* w4_rsc_61_0     [130] */ , 
    ACTIVE /* w4_rsc_62_0     [131] */ , 
    ACTIVE /* w4_rsc_63_0     [132] */ , 
    ACTIVE /* b4_rsc     [133] */ , 
    ACTIVE /* w6_rsc_0_0     [134] */ , 
    ACTIVE /* w6_rsc_1_0     [135] */ , 
    ACTIVE /* w6_rsc_2_0     [136] */ , 
    ACTIVE /* w6_rsc_3_0     [137] */ , 
    ACTIVE /* w6_rsc_4_0     [138] */ , 
    ACTIVE /* w6_rsc_5_0     [139] */ , 
    ACTIVE /* w6_rsc_6_0     [140] */ , 
    ACTIVE /* w6_rsc_7_0     [141] */ , 
    ACTIVE /* w6_rsc_8_0     [142] */ , 
    ACTIVE /* w6_rsc_9_0     [143] */ , 
    ACTIVE /* b6_rsc     [144] */   };

  // ****************************************************************************
  // FUNCTION: new()
  // This is the standard system verilog constructor.  All components are 
  // constructed in the build_phase to allow factory overriding.
  //
  function new( string name = "", uvm_component parent = null );
     super.new( name ,parent );
  endfunction



  // ****************************************************************************
  // FUNCTION: build_phase()
  // The construction of the configuration and environment classes is done in
  // the build_phase of uvmf_test_base.  Once the configuraton and environment
  // classes are built then the initialize call is made to perform the
  // following: 
  //     Monitor and driver BFM virtual interface handle passing into agents
  //     Set the active/passive state for each agent
  // Once this build_phase completes, the build_phase of the environment is
  // executed which builds the agents.
  //
  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    configuration.initialize(BLOCK, "uvm_test_top.environment", interface_names, null, interface_activities);
  endfunction

endclass
